magic
tech sky130A
magscale 1 2
timestamp 1717891028
<< error_s >>
rect -12840 -50258 -12758 -49938
rect -12520 -50258 -12438 -49938
rect -11040 -50258 -10958 -49938
rect -10720 -50258 -10638 -49938
rect -9240 -50258 -9158 -49938
rect -8920 -50258 -8838 -49938
rect -7440 -50258 -7358 -49938
rect -7120 -50258 -7038 -49938
rect -5640 -50258 -5558 -49938
rect -5320 -50258 -5238 -49938
rect -3840 -50258 -3758 -49938
rect -3520 -50258 -3438 -49938
rect -2040 -50258 -1958 -49938
rect -1720 -50258 -1638 -49938
rect -240 -50258 -158 -49938
rect 80 -50258 162 -49938
rect 1560 -50258 1642 -49938
rect 1880 -50258 1962 -49938
rect -12840 -52756 -12758 -52436
rect -12520 -52756 -12438 -52436
rect -11040 -52756 -10958 -52436
rect -10720 -52756 -10638 -52436
rect -9240 -52756 -9158 -52436
rect -8920 -52756 -8838 -52436
rect -7440 -52756 -7358 -52436
rect -7120 -52756 -7038 -52436
rect -5640 -52756 -5558 -52436
rect -5320 -52756 -5238 -52436
rect -3840 -52756 -3758 -52436
rect -3520 -52756 -3438 -52436
rect -2040 -52756 -1958 -52436
rect -1720 -52756 -1638 -52436
rect -240 -52756 -158 -52436
rect 80 -52756 162 -52436
rect 1560 -52756 1642 -52436
rect 1880 -52756 1962 -52436
rect -12840 -55254 -12758 -54934
rect -12520 -55254 -12438 -54934
rect -11040 -55254 -10958 -54934
rect -10720 -55254 -10638 -54934
rect -9240 -55254 -9158 -54934
rect -8920 -55254 -8838 -54934
rect -7440 -55254 -7358 -54934
rect -7120 -55254 -7038 -54934
rect -5640 -55254 -5558 -54934
rect -5320 -55254 -5238 -54934
rect -3840 -55254 -3758 -54934
rect -3520 -55254 -3438 -54934
rect -2040 -55254 -1958 -54934
rect -1720 -55254 -1638 -54934
rect -240 -55254 -158 -54934
rect 80 -55254 162 -54934
rect 1560 -55254 1642 -54934
rect 1880 -55254 1962 -54934
rect -12840 -57752 -12758 -57432
rect -12520 -57752 -12438 -57432
rect -11040 -57752 -10958 -57432
rect -10720 -57752 -10638 -57432
rect -9240 -57752 -9158 -57432
rect -8920 -57752 -8838 -57432
rect -7440 -57752 -7358 -57432
rect -7120 -57752 -7038 -57432
rect -5640 -57752 -5558 -57432
rect -5320 -57752 -5238 -57432
rect -3840 -57752 -3758 -57432
rect -3520 -57752 -3438 -57432
rect -2040 -57752 -1958 -57432
rect -1720 -57752 -1638 -57432
rect -240 -57752 -158 -57432
rect 80 -57752 162 -57432
rect 1560 -57752 1642 -57432
rect 1880 -57752 1962 -57432
rect -12840 -60250 -12758 -59930
rect -12520 -60250 -12438 -59930
rect -11040 -60250 -10958 -59930
rect -10720 -60250 -10638 -59930
rect -9240 -60250 -9158 -59930
rect -8920 -60250 -8838 -59930
rect -7440 -60250 -7358 -59930
rect -7120 -60250 -7038 -59930
rect -5640 -60250 -5558 -59930
rect -5320 -60250 -5238 -59930
rect -3840 -60250 -3758 -59930
rect -3520 -60250 -3438 -59930
rect -2040 -60250 -1958 -59930
rect -1720 -60250 -1638 -59930
rect -240 -60250 -158 -59930
rect 80 -60250 162 -59930
rect 1560 -60250 1642 -59930
rect 1880 -60250 1962 -59930
rect -12840 -62748 -12758 -62428
rect -12520 -62748 -12438 -62428
rect -11040 -62748 -10958 -62428
rect -10720 -62748 -10638 -62428
rect -9240 -62748 -9158 -62428
rect -8920 -62748 -8838 -62428
rect -7440 -62748 -7358 -62428
rect -7120 -62748 -7038 -62428
rect -5640 -62748 -5558 -62428
rect -5320 -62748 -5238 -62428
rect -3840 -62748 -3758 -62428
rect -3520 -62748 -3438 -62428
rect -2040 -62748 -1958 -62428
rect -1720 -62748 -1638 -62428
rect -240 -62748 -158 -62428
rect 80 -62748 162 -62428
rect 1560 -62748 1642 -62428
rect 1880 -62748 1962 -62428
rect -12840 -65246 -12758 -64926
rect -12520 -65246 -12438 -64926
rect -11040 -65246 -10958 -64926
rect -10720 -65246 -10638 -64926
rect -9240 -65246 -9158 -64926
rect -8920 -65246 -8838 -64926
rect -7440 -65246 -7358 -64926
rect -7120 -65246 -7038 -64926
rect -5640 -65246 -5558 -64926
rect -5320 -65246 -5238 -64926
rect -3840 -65246 -3758 -64926
rect -3520 -65246 -3438 -64926
rect -2040 -65246 -1958 -64926
rect -1720 -65246 -1638 -64926
rect -240 -65246 -158 -64926
rect 80 -65246 162 -64926
rect 1560 -65246 1642 -64926
rect 1880 -65246 1962 -64926
rect -12840 -67744 -12758 -67424
rect -12520 -67744 -12438 -67424
rect -11040 -67744 -10958 -67424
rect -10720 -67744 -10638 -67424
rect -9240 -67744 -9158 -67424
rect -8920 -67744 -8838 -67424
rect -7440 -67744 -7358 -67424
rect -7120 -67744 -7038 -67424
rect -5640 -67744 -5558 -67424
rect -5320 -67744 -5238 -67424
rect -3840 -67744 -3758 -67424
rect -3520 -67744 -3438 -67424
rect -2040 -67744 -1958 -67424
rect -1720 -67744 -1638 -67424
rect -240 -67744 -158 -67424
rect 80 -67744 162 -67424
rect 1560 -67744 1642 -67424
rect 1880 -67744 1962 -67424
rect -12840 -70242 -12758 -69922
rect -12520 -70242 -12438 -69922
rect -11040 -70242 -10958 -69922
rect -10720 -70242 -10638 -69922
rect -9240 -70242 -9158 -69922
rect -8920 -70242 -8838 -69922
rect -7440 -70242 -7358 -69922
rect -7120 -70242 -7038 -69922
rect -5640 -70242 -5558 -69922
rect -5320 -70242 -5238 -69922
rect -3840 -70242 -3758 -69922
rect -3520 -70242 -3438 -69922
rect -2040 -70242 -1958 -69922
rect -1720 -70242 -1638 -69922
rect -240 -70242 -158 -69922
rect 80 -70242 162 -69922
rect 1560 -70242 1642 -69922
rect 1880 -70242 1962 -69922
<< metal1 >>
rect -15196 -60838 -14996 -60638
rect -15196 -61238 -14996 -61038
rect -15196 -61638 -14996 -61438
rect -15196 -62038 -14996 -61838
rect -15196 -62438 -14996 -62238
rect -15196 -62838 -14996 -62638
rect -15196 -63238 -14996 -63038
use sky130_fd_pr__cap_mim_m3_1_4ABMPW  sky130_fd_pr__cap_mim_m3_1_4ABMPW_0 paramcells
timestamp 1717890828
transform 0 1 -5799 -1 0 -59472
box -8934 -8480 12822 9200
use sky130_fd_pr__cap_mim_m3_2_4ABMPW  XC4 paramcells
timestamp 1717881426
transform 0 -1 -5439 1 0 -61001
box -11041 -8881 11063 8881
<< labels >>
flabel metal1 -15196 -60838 -14996 -60638 0 FreeSans 256 0 0 0 D8
port 0 nsew
flabel metal1 -15196 -61238 -14996 -61038 0 FreeSans 256 0 0 0 D5
port 1 nsew
flabel metal1 -15196 -61638 -14996 -61438 0 FreeSans 256 0 0 0 D9
port 2 nsew
flabel metal1 -15196 -62038 -14996 -61838 0 FreeSans 256 0 0 0 VP2
port 3 nsew
flabel metal1 -15196 -62438 -14996 -62238 0 FreeSans 256 0 0 0 D6
port 4 nsew
flabel metal1 -15196 -62838 -14996 -62638 0 FreeSans 256 0 0 0 VSS
port 5 nsew
flabel metal1 -15196 -63238 -14996 -63038 0 FreeSans 256 0 0 0 D7
port 6 nsew
<< end >>
