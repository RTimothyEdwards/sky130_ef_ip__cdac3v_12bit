magic
tech sky130A
magscale 1 2
timestamp 1717890828
<< error_s >>
rect -10511 -19078 -10429 -18758
rect -10191 -19078 -10109 -18758
rect -8711 -19078 -8629 -18758
rect -8391 -19078 -8309 -18758
rect -6911 -19078 -6829 -18758
rect -6591 -19078 -6509 -18758
rect -5111 -19078 -5029 -18758
rect -4791 -19078 -4709 -18758
rect -3311 -19078 -3229 -18758
rect -2991 -19078 -2909 -18758
rect -1511 -19078 -1429 -18758
rect -1191 -19078 -1109 -18758
rect 289 -19078 371 -18758
rect 609 -19078 691 -18758
rect 2089 -19078 2171 -18758
rect 2409 -19078 2491 -18758
rect 3889 -19078 3971 -18758
rect 4209 -19078 4291 -18758
rect -10511 -21576 -10429 -21256
rect -10191 -21576 -10109 -21256
rect -8711 -21576 -8629 -21256
rect -8391 -21576 -8309 -21256
rect -6911 -21576 -6829 -21256
rect -6591 -21576 -6509 -21256
rect -5111 -21576 -5029 -21256
rect -4791 -21576 -4709 -21256
rect -3311 -21576 -3229 -21256
rect -2991 -21576 -2909 -21256
rect -1511 -21576 -1429 -21256
rect -1191 -21576 -1109 -21256
rect 289 -21576 371 -21256
rect 609 -21576 691 -21256
rect 2089 -21576 2171 -21256
rect 2409 -21576 2491 -21256
rect 3889 -21576 3971 -21256
rect 4209 -21576 4291 -21256
rect -10511 -24074 -10429 -23754
rect -10191 -24074 -10109 -23754
rect -8711 -24074 -8629 -23754
rect -8391 -24074 -8309 -23754
rect -6911 -24074 -6829 -23754
rect -6591 -24074 -6509 -23754
rect -5111 -24074 -5029 -23754
rect -4791 -24074 -4709 -23754
rect -3311 -24074 -3229 -23754
rect -2991 -24074 -2909 -23754
rect -1511 -24074 -1429 -23754
rect -1191 -24074 -1109 -23754
rect 289 -24074 371 -23754
rect 609 -24074 691 -23754
rect 2089 -24074 2171 -23754
rect 2409 -24074 2491 -23754
rect 3889 -24074 3971 -23754
rect 4209 -24074 4291 -23754
rect -10511 -26572 -10429 -26252
rect -10191 -26572 -10109 -26252
rect -8711 -26572 -8629 -26252
rect -8391 -26572 -8309 -26252
rect -6911 -26572 -6829 -26252
rect -6591 -26572 -6509 -26252
rect -5111 -26572 -5029 -26252
rect -4791 -26572 -4709 -26252
rect -3311 -26572 -3229 -26252
rect -2991 -26572 -2909 -26252
rect -1511 -26572 -1429 -26252
rect -1191 -26572 -1109 -26252
rect 289 -26572 371 -26252
rect 609 -26572 691 -26252
rect 2089 -26572 2171 -26252
rect 2409 -26572 2491 -26252
rect 3889 -26572 3971 -26252
rect 4209 -26572 4291 -26252
rect -10511 -29070 -10429 -28750
rect -10191 -29070 -10109 -28750
rect -8711 -29070 -8629 -28750
rect -8391 -29070 -8309 -28750
rect -6911 -29070 -6829 -28750
rect -6591 -29070 -6509 -28750
rect -5111 -29070 -5029 -28750
rect -4791 -29070 -4709 -28750
rect -3311 -29070 -3229 -28750
rect -2991 -29070 -2909 -28750
rect -1511 -29070 -1429 -28750
rect -1191 -29070 -1109 -28750
rect 289 -29070 371 -28750
rect 609 -29070 691 -28750
rect 2089 -29070 2171 -28750
rect 2409 -29070 2491 -28750
rect 3889 -29070 3971 -28750
rect 4209 -29070 4291 -28750
rect -10511 -31568 -10429 -31248
rect -10191 -31568 -10109 -31248
rect -8711 -31568 -8629 -31248
rect -8391 -31568 -8309 -31248
rect -6911 -31568 -6829 -31248
rect -6591 -31568 -6509 -31248
rect -5111 -31568 -5029 -31248
rect -4791 -31568 -4709 -31248
rect -3311 -31568 -3229 -31248
rect -2991 -31568 -2909 -31248
rect -1511 -31568 -1429 -31248
rect -1191 -31568 -1109 -31248
rect 289 -31568 371 -31248
rect 609 -31568 691 -31248
rect 2089 -31568 2171 -31248
rect 2409 -31568 2491 -31248
rect 3889 -31568 3971 -31248
rect 4209 -31568 4291 -31248
rect -10511 -34066 -10429 -33746
rect -10191 -34066 -10109 -33746
rect -8711 -34066 -8629 -33746
rect -8391 -34066 -8309 -33746
rect -6911 -34066 -6829 -33746
rect -6591 -34066 -6509 -33746
rect -5111 -34066 -5029 -33746
rect -4791 -34066 -4709 -33746
rect -3311 -34066 -3229 -33746
rect -2991 -34066 -2909 -33746
rect -1511 -34066 -1429 -33746
rect -1191 -34066 -1109 -33746
rect 289 -34066 371 -33746
rect 609 -34066 691 -33746
rect 2089 -34066 2171 -33746
rect 2409 -34066 2491 -33746
rect 3889 -34066 3971 -33746
rect 4209 -34066 4291 -33746
rect -10511 -36564 -10429 -36244
rect -10191 -36564 -10109 -36244
rect -8711 -36564 -8629 -36244
rect -8391 -36564 -8309 -36244
rect -6911 -36564 -6829 -36244
rect -6591 -36564 -6509 -36244
rect -5111 -36564 -5029 -36244
rect -4791 -36564 -4709 -36244
rect -3311 -36564 -3229 -36244
rect -2991 -36564 -2909 -36244
rect -1511 -36564 -1429 -36244
rect -1191 -36564 -1109 -36244
rect 289 -36564 371 -36244
rect 609 -36564 691 -36244
rect 2089 -36564 2171 -36244
rect 2409 -36564 2491 -36244
rect 3889 -36564 3971 -36244
rect 4209 -36564 4291 -36244
rect -10511 -39062 -10429 -38742
rect -10191 -39062 -10109 -38742
rect -8711 -39062 -8629 -38742
rect -8391 -39062 -8309 -38742
rect -6911 -39062 -6829 -38742
rect -6591 -39062 -6509 -38742
rect -5111 -39062 -5029 -38742
rect -4791 -39062 -4709 -38742
rect -3311 -39062 -3229 -38742
rect -2991 -39062 -2909 -38742
rect -1511 -39062 -1429 -38742
rect -1191 -39062 -1109 -38742
rect 289 -39062 371 -38742
rect 609 -39062 691 -38742
rect 2089 -39062 2171 -38742
rect 2409 -39062 2491 -38742
rect 3889 -39062 3971 -38742
rect 4209 -39062 4291 -38742
<< metal1 >>
rect -14578 -29154 -14378 -28954
rect -14578 -29554 -14378 -29354
rect -14578 -29954 -14378 -29754
rect -14578 -30354 -14378 -30154
rect -14578 -30754 -14378 -30554
rect -14578 -31154 -14378 -30954
rect -14578 -31554 -14378 -31354
use sky130_fd_pr__cap_mim_m3_2_4ABMPW  sky130_fd_pr__cap_mim_m3_2_4ABMPW_0 paramcells
timestamp 1717881426
transform 0 -1 -3110 1 0 -29821
box -11041 -8881 11063 8881
use sky130_fd_pr__cap_mim_m3_1_4ABMPW  XC6 paramcells
timestamp 1717890828
transform 0 1 -3470 -1 0 -28292
box -8934 -8480 12822 9200
<< labels >>
flabel metal1 -14578 -29154 -14378 -28954 0 FreeSans 256 0 0 0 VP1
port 0 nsew
flabel metal1 -14578 -29554 -14378 -29354 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 -14578 -29954 -14378 -29754 0 FreeSans 256 0 0 0 D0
port 2 nsew
flabel metal1 -14578 -30354 -14378 -30154 0 FreeSans 256 0 0 0 D1
port 3 nsew
flabel metal1 -14578 -30754 -14378 -30554 0 FreeSans 256 0 0 0 D2
port 4 nsew
flabel metal1 -14578 -31154 -14378 -30954 0 FreeSans 256 0 0 0 D3
port 5 nsew
flabel metal1 -14578 -31554 -14378 -31354 0 FreeSans 256 0 0 0 D4
port 6 nsew
<< end >>
