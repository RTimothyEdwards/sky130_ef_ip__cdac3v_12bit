magic
tech sky130A
magscale 1 2
timestamp 1722437419
<< metal1 >>
rect 5959 27041 6159 27241
rect 12963 27041 13163 27241
rect 19967 27041 20167 27241
rect 33975 27041 34175 27241
rect 40979 27041 41179 27241
rect 47983 27041 48183 27241
rect 5959 -8994 6159 -8794
rect 12963 -8994 13163 -8794
rect 19967 -8994 20167 -8794
rect 33975 -8994 34175 -8794
rect 40979 -8994 41179 -8794
rect 47983 -8994 48183 -8794
<< via2 >>
rect 7209 23783 7399 23933
rect 14213 23783 14403 23933
rect 21217 23783 21407 23933
rect 35225 23783 35415 23933
rect 42229 23783 42419 23933
rect 49233 23783 49423 23933
rect 1790 23485 1980 23635
rect 8794 23485 8984 23635
rect 15798 23485 15988 23635
rect 29806 23485 29996 23635
rect 36810 23485 37000 23635
rect 43814 23485 44004 23635
rect 1790 -5387 1980 -5237
rect 8794 -5387 8984 -5237
rect 15798 -5387 15988 -5237
rect 29806 -5387 29996 -5237
rect 36810 -5387 37000 -5237
rect 43814 -5387 44004 -5237
rect 7209 -5685 7399 -5535
rect 14213 -5685 14403 -5535
rect 21217 -5685 21407 -5535
rect 35225 -5685 35415 -5535
rect 42229 -5685 42419 -5535
rect 49233 -5685 49423 -5535
<< metal3 >>
rect 22121 25897 29057 26297
rect 50155 25897 51588 26297
rect 22121 25297 29057 25697
rect 50155 25297 50967 25697
rect 320 24697 1082 25097
rect 22121 24697 29057 25097
rect 320 -6450 720 24697
rect 889 -5850 1289 24497
rect 22121 24097 29057 24497
rect 1451 23933 50352 23946
rect 1451 23783 7209 23933
rect 7399 23783 14213 23933
rect 14403 23783 21217 23933
rect 21407 23783 35225 23933
rect 35415 23783 42229 23933
rect 42419 23783 49233 23933
rect 49423 23783 50352 23933
rect 1451 23766 50352 23783
rect 1451 23635 50052 23646
rect 1451 23485 1790 23635
rect 1980 23485 8794 23635
rect 8984 23485 15798 23635
rect 15988 23485 29806 23635
rect 29996 23485 36810 23635
rect 37000 23485 43814 23635
rect 44004 23485 50052 23635
rect 1451 23466 50052 23485
rect 26832 23316 26977 23466
rect 5891 23116 6091 23316
rect 12895 23116 13095 23316
rect 19899 23116 20099 23316
rect 22179 23120 29073 23316
rect 33907 23116 34107 23316
rect 40911 23116 41111 23316
rect 47915 23116 48115 23316
rect 49872 8764 50052 23466
rect 50172 9164 50352 23766
rect 50131 8964 50352 9164
rect 49851 8564 50052 8764
rect 5891 -5069 6091 -4869
rect 12895 -5069 13095 -4869
rect 19899 -5069 20099 -4869
rect 33907 -5069 34107 -4869
rect 40911 -5069 41111 -4869
rect 47915 -5069 48115 -4869
rect 49872 -5221 50052 8564
rect 1451 -5237 50052 -5221
rect 1451 -5387 1790 -5237
rect 1980 -5387 8794 -5237
rect 8984 -5387 15798 -5237
rect 15988 -5387 29806 -5237
rect 29996 -5387 36810 -5237
rect 37000 -5387 43814 -5237
rect 44004 -5387 50052 -5237
rect 1451 -5401 50052 -5387
rect 50172 -5521 50352 8964
rect 1451 -5535 50352 -5521
rect 1451 -5685 7209 -5535
rect 7399 -5685 14213 -5535
rect 14403 -5685 21217 -5535
rect 21407 -5685 35225 -5535
rect 35415 -5685 42229 -5535
rect 42419 -5685 49233 -5535
rect 49423 -5685 50352 -5535
rect 1451 -5701 50352 -5685
rect 889 -6250 1301 -5850
rect 22123 -6250 29049 -5850
rect 50154 -6250 50436 -5850
rect 320 -6850 1301 -6450
rect 22123 -6850 29049 -6450
rect 50154 -6850 50436 -6450
rect 50567 -7050 50967 25297
rect 22142 -7450 29058 -7050
rect 50074 -7450 50967 -7050
rect 51188 -7650 51588 25897
rect 22142 -8050 29058 -7650
rect 50074 -8050 51588 -7650
use EF_AMUX21x  EF_AMUX21x_0
timestamp 1722435879
transform 0 -1 13438 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  EF_AMUX21x_1
timestamp 1722435879
transform 0 -1 6434 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  x1
timestamp 1722435879
transform 0 -1 27446 -1 0 27907
box 656 -8770 5084 -1560
use EF_AMUX21x  x2
timestamp 1722435879
transform 0 -1 41454 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  x3
timestamp 1722435879
transform 0 -1 13438 -1 0 27907
box 656 -8770 5084 -1560
use EF_AMUX21x  x4
timestamp 1722435879
transform 0 -1 6434 -1 0 27907
box 656 -8770 5084 -1560
use EF_AMUX21x  x5
timestamp 1722435879
transform 0 -1 34450 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  x8
timestamp 1722435879
transform 0 -1 27446 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  x9
timestamp 1722435879
transform 0 -1 -570 1 0 -9660
box 656 -8770 5084 -1560
use EF_AMUX21x  x10
timestamp 1722435879
transform 0 -1 41454 -1 0 27907
box 656 -8770 5084 -1560
use EF_AMUX21x  x11
timestamp 1722435879
transform 0 -1 34450 -1 0 27907
box 656 -8770 5084 -1560
use EF_AMUX21x  x12
timestamp 1722435879
transform 0 -1 -570 -1 0 27907
box 656 -8770 5084 -1560
<< labels >>
flabel metal1 5959 -8994 6159 -8794 0 FreeSans 256 90 0 0 SELD11
port 30 nsew
flabel metal1 12963 -8994 13163 -8794 0 FreeSans 256 90 0 0 SELD7
port 14 nsew
flabel metal1 19967 -8994 20167 -8794 0 FreeSans 256 90 0 0 SELD9
port 11 nsew
flabel metal1 33975 -8994 34175 -8794 0 FreeSans 256 90 0 0 SELD2
port 1 nsew
flabel metal1 40979 -8994 41179 -8794 0 FreeSans 256 90 0 0 SELD0
port 4 nsew
flabel metal1 47983 -8994 48183 -8794 0 FreeSans 256 90 0 0 SELD4
port 7 nsew
flabel metal3 5891 -5069 6091 -4869 0 FreeSans 256 90 0 0 D11
port 28 nsew
flabel metal3 12895 -5069 13095 -4869 0 FreeSans 256 90 0 0 D7
port 18 nsew
flabel metal3 19899 -5069 20099 -4869 0 FreeSans 256 90 0 0 D9
port 15 nsew
flabel metal3 33907 -5069 34107 -4869 0 FreeSans 256 90 0 0 D2
port 0 nsew
flabel metal3 40911 -5069 41111 -4869 0 FreeSans 256 90 0 0 D0
port 5 nsew
flabel metal3 47915 -5069 48115 -4869 0 FreeSans 256 90 0 0 D4
port 10 nsew
flabel metal3 50235 -6747 50435 -6547 0 FreeSans 256 180 0 0 DVDD
port 21 nsew
flabel metal3 50237 -7341 50437 -7141 0 FreeSans 256 180 0 0 VSS
port 26 nsew
flabel metal3 50237 -7934 50437 -7734 0 FreeSans 256 180 0 0 VDD
port 20 nsew
flabel metal3 50233 -6176 50433 -5976 0 FreeSans 256 180 0 0 DVSS
port 22 nsew
flabel metal1 47983 27041 48183 27241 0 FreeSans 256 90 0 0 SELD5
port 9 nsew
flabel metal1 40979 27041 41179 27241 0 FreeSans 256 90 0 0 SELD1
port 6 nsew
flabel metal1 33975 27041 34175 27241 0 FreeSans 256 90 0 0 SELD3
port 3 nsew
flabel metal1 19967 27041 20167 27241 0 FreeSans 256 90 0 0 SELD8
port 12 nsew
flabel metal1 5959 27041 6159 27241 0 FreeSans 256 90 0 0 SELD10
port 29 nsew
flabel metal1 12963 27041 13163 27241 0 FreeSans 256 90 0 0 SELD6
port 16 nsew
flabel metal3 5891 23116 6091 23316 0 FreeSans 256 90 0 0 D10
port 27 nsew
flabel metal3 12895 23116 13095 23316 0 FreeSans 256 90 0 0 D6
port 19 nsew
flabel metal3 19899 23116 20099 23316 0 FreeSans 256 90 0 0 D8
port 17 nsew
flabel metal3 33907 23116 34107 23316 0 FreeSans 256 90 0 0 D3
port 2 nsew
flabel metal3 40911 23116 41111 23316 0 FreeSans 256 90 0 0 D1
port 8 nsew
flabel metal3 47915 23116 48115 23316 0 FreeSans 256 90 0 0 D5
port 13 nsew
flabel metal3 50131 8964 50331 9164 0 FreeSans 256 180 0 0 VH
port 24 nsew
flabel metal3 49851 8564 50051 8764 0 FreeSans 256 180 0 0 VL
port 25 nsew
<< end >>
