magic
tech sky130A
magscale 1 2
timestamp 1717881426
<< error_p >>
rect -9241 7319 -8921 7401
rect -6743 7319 -6423 7401
rect -4245 7319 -3925 7401
rect -1747 7319 -1427 7401
rect 751 7319 1071 7401
rect 3249 7319 3569 7401
rect 5747 7319 6067 7401
rect 8245 7319 8565 7401
rect 10743 7319 11063 7401
rect -9241 6999 -8921 7081
rect -6743 6999 -6423 7081
rect -4245 6999 -3925 7081
rect -1747 6999 -1427 7081
rect 751 6999 1071 7081
rect 3249 6999 3569 7081
rect 5747 6999 6067 7081
rect 8245 6999 8565 7081
rect 10743 6999 11063 7081
rect -9241 5519 -8921 5601
rect -6743 5519 -6423 5601
rect -4245 5519 -3925 5601
rect -1747 5519 -1427 5601
rect 751 5519 1071 5601
rect 3249 5519 3569 5601
rect 5747 5519 6067 5601
rect 8245 5519 8565 5601
rect 10743 5519 11063 5601
rect -9241 5199 -8921 5281
rect -6743 5199 -6423 5281
rect -4245 5199 -3925 5281
rect -1747 5199 -1427 5281
rect 751 5199 1071 5281
rect 3249 5199 3569 5281
rect 5747 5199 6067 5281
rect 8245 5199 8565 5281
rect 10743 5199 11063 5281
rect -9241 3719 -8921 3801
rect -6743 3719 -6423 3801
rect -4245 3719 -3925 3801
rect -1747 3719 -1427 3801
rect 751 3719 1071 3801
rect 3249 3719 3569 3801
rect 5747 3719 6067 3801
rect 8245 3719 8565 3801
rect 10743 3719 11063 3801
rect -9241 3399 -8921 3481
rect -6743 3399 -6423 3481
rect -4245 3399 -3925 3481
rect -1747 3399 -1427 3481
rect 751 3399 1071 3481
rect 3249 3399 3569 3481
rect 5747 3399 6067 3481
rect 8245 3399 8565 3481
rect 10743 3399 11063 3481
rect -9241 1919 -8921 2001
rect -6743 1919 -6423 2001
rect -4245 1919 -3925 2001
rect -1747 1919 -1427 2001
rect 751 1919 1071 2001
rect 3249 1919 3569 2001
rect 5747 1919 6067 2001
rect 8245 1919 8565 2001
rect 10743 1919 11063 2001
rect -9241 1599 -8921 1681
rect -6743 1599 -6423 1681
rect -4245 1599 -3925 1681
rect -1747 1599 -1427 1681
rect 751 1599 1071 1681
rect 3249 1599 3569 1681
rect 5747 1599 6067 1681
rect 8245 1599 8565 1681
rect 10743 1599 11063 1681
rect -9241 119 -8921 201
rect -6743 119 -6423 201
rect -4245 119 -3925 201
rect -1747 119 -1427 201
rect 751 119 1071 201
rect 3249 119 3569 201
rect 5747 119 6067 201
rect 8245 119 8565 201
rect 10743 119 11063 201
rect -9241 -201 -8921 -119
rect -6743 -201 -6423 -119
rect -4245 -201 -3925 -119
rect -1747 -201 -1427 -119
rect 751 -201 1071 -119
rect 3249 -201 3569 -119
rect 5747 -201 6067 -119
rect 8245 -201 8565 -119
rect 10743 -201 11063 -119
rect -9241 -1681 -8921 -1599
rect -6743 -1681 -6423 -1599
rect -4245 -1681 -3925 -1599
rect -1747 -1681 -1427 -1599
rect 751 -1681 1071 -1599
rect 3249 -1681 3569 -1599
rect 5747 -1681 6067 -1599
rect 8245 -1681 8565 -1599
rect 10743 -1681 11063 -1599
rect -9241 -2001 -8921 -1919
rect -6743 -2001 -6423 -1919
rect -4245 -2001 -3925 -1919
rect -1747 -2001 -1427 -1919
rect 751 -2001 1071 -1919
rect 3249 -2001 3569 -1919
rect 5747 -2001 6067 -1919
rect 8245 -2001 8565 -1919
rect 10743 -2001 11063 -1919
rect -9241 -3481 -8921 -3399
rect -6743 -3481 -6423 -3399
rect -4245 -3481 -3925 -3399
rect -1747 -3481 -1427 -3399
rect 751 -3481 1071 -3399
rect 3249 -3481 3569 -3399
rect 5747 -3481 6067 -3399
rect 8245 -3481 8565 -3399
rect 10743 -3481 11063 -3399
rect -9241 -3801 -8921 -3719
rect -6743 -3801 -6423 -3719
rect -4245 -3801 -3925 -3719
rect -1747 -3801 -1427 -3719
rect 751 -3801 1071 -3719
rect 3249 -3801 3569 -3719
rect 5747 -3801 6067 -3719
rect 8245 -3801 8565 -3719
rect 10743 -3801 11063 -3719
rect -9241 -5281 -8921 -5199
rect -6743 -5281 -6423 -5199
rect -4245 -5281 -3925 -5199
rect -1747 -5281 -1427 -5199
rect 751 -5281 1071 -5199
rect 3249 -5281 3569 -5199
rect 5747 -5281 6067 -5199
rect 8245 -5281 8565 -5199
rect 10743 -5281 11063 -5199
rect -9241 -5601 -8921 -5519
rect -6743 -5601 -6423 -5519
rect -4245 -5601 -3925 -5519
rect -1747 -5601 -1427 -5519
rect 751 -5601 1071 -5519
rect 3249 -5601 3569 -5519
rect 5747 -5601 6067 -5519
rect 8245 -5601 8565 -5519
rect 10743 -5601 11063 -5519
rect -9241 -7081 -8921 -6999
rect -6743 -7081 -6423 -6999
rect -4245 -7081 -3925 -6999
rect -1747 -7081 -1427 -6999
rect 751 -7081 1071 -6999
rect 3249 -7081 3569 -6999
rect 5747 -7081 6067 -6999
rect 8245 -7081 8565 -6999
rect 10743 -7081 11063 -6999
rect -9241 -7401 -8921 -7319
rect -6743 -7401 -6423 -7319
rect -4245 -7401 -3925 -7319
rect -1747 -7401 -1427 -7319
rect 751 -7401 1071 -7319
rect 3249 -7401 3569 -7319
rect 5747 -7401 6067 -7319
rect 8245 -7401 8565 -7319
rect 10743 -7401 11063 -7319
<< metal4 >>
rect -11041 8839 -8943 8880
rect -11041 7361 -9199 8839
rect -8963 7361 -8943 8839
rect -11041 7320 -8943 7361
rect -8543 8839 -6445 8880
rect -8543 7361 -6701 8839
rect -6465 7361 -6445 8839
rect -8543 7320 -6445 7361
rect -6045 8839 -3947 8880
rect -6045 7361 -4203 8839
rect -3967 7361 -3947 8839
rect -6045 7320 -3947 7361
rect -3547 8839 -1449 8880
rect -3547 7361 -1705 8839
rect -1469 7361 -1449 8839
rect -3547 7320 -1449 7361
rect -1049 8839 1049 8880
rect -1049 7361 793 8839
rect 1029 7361 1049 8839
rect -1049 7320 1049 7361
rect 1449 8839 3547 8880
rect 1449 7361 3291 8839
rect 3527 7361 3547 8839
rect 1449 7320 3547 7361
rect 3947 8839 6045 8880
rect 3947 7361 5789 8839
rect 6025 7361 6045 8839
rect 3947 7320 6045 7361
rect 6445 8839 8543 8880
rect 6445 7361 8287 8839
rect 8523 7361 8543 8839
rect 6445 7320 8543 7361
rect 8943 8839 11041 8880
rect 8943 7361 10785 8839
rect 11021 7361 11041 8839
rect 8943 7320 11041 7361
rect -11041 7039 -8943 7080
rect -11041 5561 -9199 7039
rect -8963 5561 -8943 7039
rect -11041 5520 -8943 5561
rect -8543 7039 -6445 7080
rect -8543 5561 -6701 7039
rect -6465 5561 -6445 7039
rect -8543 5520 -6445 5561
rect -6045 7039 -3947 7080
rect -6045 5561 -4203 7039
rect -3967 5561 -3947 7039
rect -6045 5520 -3947 5561
rect -3547 7039 -1449 7080
rect -3547 5561 -1705 7039
rect -1469 5561 -1449 7039
rect -3547 5520 -1449 5561
rect -1049 7039 1049 7080
rect -1049 5561 793 7039
rect 1029 5561 1049 7039
rect -1049 5520 1049 5561
rect 1449 7039 3547 7080
rect 1449 5561 3291 7039
rect 3527 5561 3547 7039
rect 1449 5520 3547 5561
rect 3947 7039 6045 7080
rect 3947 5561 5789 7039
rect 6025 5561 6045 7039
rect 3947 5520 6045 5561
rect 6445 7039 8543 7080
rect 6445 5561 8287 7039
rect 8523 5561 8543 7039
rect 6445 5520 8543 5561
rect 8943 7039 11041 7080
rect 8943 5561 10785 7039
rect 11021 5561 11041 7039
rect 8943 5520 11041 5561
rect -11041 5239 -8943 5280
rect -11041 3761 -9199 5239
rect -8963 3761 -8943 5239
rect -11041 3720 -8943 3761
rect -8543 5239 -6445 5280
rect -8543 3761 -6701 5239
rect -6465 3761 -6445 5239
rect -8543 3720 -6445 3761
rect -6045 5239 -3947 5280
rect -6045 3761 -4203 5239
rect -3967 3761 -3947 5239
rect -6045 3720 -3947 3761
rect -3547 5239 -1449 5280
rect -3547 3761 -1705 5239
rect -1469 3761 -1449 5239
rect -3547 3720 -1449 3761
rect -1049 5239 1049 5280
rect -1049 3761 793 5239
rect 1029 3761 1049 5239
rect -1049 3720 1049 3761
rect 1449 5239 3547 5280
rect 1449 3761 3291 5239
rect 3527 3761 3547 5239
rect 1449 3720 3547 3761
rect 3947 5239 6045 5280
rect 3947 3761 5789 5239
rect 6025 3761 6045 5239
rect 3947 3720 6045 3761
rect 6445 5239 8543 5280
rect 6445 3761 8287 5239
rect 8523 3761 8543 5239
rect 6445 3720 8543 3761
rect 8943 5239 11041 5280
rect 8943 3761 10785 5239
rect 11021 3761 11041 5239
rect 8943 3720 11041 3761
rect -11041 3439 -8943 3480
rect -11041 1961 -9199 3439
rect -8963 1961 -8943 3439
rect -11041 1920 -8943 1961
rect -8543 3439 -6445 3480
rect -8543 1961 -6701 3439
rect -6465 1961 -6445 3439
rect -8543 1920 -6445 1961
rect -6045 3439 -3947 3480
rect -6045 1961 -4203 3439
rect -3967 1961 -3947 3439
rect -6045 1920 -3947 1961
rect -3547 3439 -1449 3480
rect -3547 1961 -1705 3439
rect -1469 1961 -1449 3439
rect -3547 1920 -1449 1961
rect -1049 3439 1049 3480
rect -1049 1961 793 3439
rect 1029 1961 1049 3439
rect -1049 1920 1049 1961
rect 1449 3439 3547 3480
rect 1449 1961 3291 3439
rect 3527 1961 3547 3439
rect 1449 1920 3547 1961
rect 3947 3439 6045 3480
rect 3947 1961 5789 3439
rect 6025 1961 6045 3439
rect 3947 1920 6045 1961
rect 6445 3439 8543 3480
rect 6445 1961 8287 3439
rect 8523 1961 8543 3439
rect 6445 1920 8543 1961
rect 8943 3439 11041 3480
rect 8943 1961 10785 3439
rect 11021 1961 11041 3439
rect 8943 1920 11041 1961
rect -11041 1639 -8943 1680
rect -11041 161 -9199 1639
rect -8963 161 -8943 1639
rect -11041 120 -8943 161
rect -8543 1639 -6445 1680
rect -8543 161 -6701 1639
rect -6465 161 -6445 1639
rect -8543 120 -6445 161
rect -6045 1639 -3947 1680
rect -6045 161 -4203 1639
rect -3967 161 -3947 1639
rect -6045 120 -3947 161
rect -3547 1639 -1449 1680
rect -3547 161 -1705 1639
rect -1469 161 -1449 1639
rect -3547 120 -1449 161
rect -1049 1639 1049 1680
rect -1049 161 793 1639
rect 1029 161 1049 1639
rect -1049 120 1049 161
rect 1449 1639 3547 1680
rect 1449 161 3291 1639
rect 3527 161 3547 1639
rect 1449 120 3547 161
rect 3947 1639 6045 1680
rect 3947 161 5789 1639
rect 6025 161 6045 1639
rect 3947 120 6045 161
rect 6445 1639 8543 1680
rect 6445 161 8287 1639
rect 8523 161 8543 1639
rect 6445 120 8543 161
rect 8943 1639 11041 1680
rect 8943 161 10785 1639
rect 11021 161 11041 1639
rect 8943 120 11041 161
rect -11041 -161 -8943 -120
rect -11041 -1639 -9199 -161
rect -8963 -1639 -8943 -161
rect -11041 -1680 -8943 -1639
rect -8543 -161 -6445 -120
rect -8543 -1639 -6701 -161
rect -6465 -1639 -6445 -161
rect -8543 -1680 -6445 -1639
rect -6045 -161 -3947 -120
rect -6045 -1639 -4203 -161
rect -3967 -1639 -3947 -161
rect -6045 -1680 -3947 -1639
rect -3547 -161 -1449 -120
rect -3547 -1639 -1705 -161
rect -1469 -1639 -1449 -161
rect -3547 -1680 -1449 -1639
rect -1049 -161 1049 -120
rect -1049 -1639 793 -161
rect 1029 -1639 1049 -161
rect -1049 -1680 1049 -1639
rect 1449 -161 3547 -120
rect 1449 -1639 3291 -161
rect 3527 -1639 3547 -161
rect 1449 -1680 3547 -1639
rect 3947 -161 6045 -120
rect 3947 -1639 5789 -161
rect 6025 -1639 6045 -161
rect 3947 -1680 6045 -1639
rect 6445 -161 8543 -120
rect 6445 -1639 8287 -161
rect 8523 -1639 8543 -161
rect 6445 -1680 8543 -1639
rect 8943 -161 11041 -120
rect 8943 -1639 10785 -161
rect 11021 -1639 11041 -161
rect 8943 -1680 11041 -1639
rect -11041 -1961 -8943 -1920
rect -11041 -3439 -9199 -1961
rect -8963 -3439 -8943 -1961
rect -11041 -3480 -8943 -3439
rect -8543 -1961 -6445 -1920
rect -8543 -3439 -6701 -1961
rect -6465 -3439 -6445 -1961
rect -8543 -3480 -6445 -3439
rect -6045 -1961 -3947 -1920
rect -6045 -3439 -4203 -1961
rect -3967 -3439 -3947 -1961
rect -6045 -3480 -3947 -3439
rect -3547 -1961 -1449 -1920
rect -3547 -3439 -1705 -1961
rect -1469 -3439 -1449 -1961
rect -3547 -3480 -1449 -3439
rect -1049 -1961 1049 -1920
rect -1049 -3439 793 -1961
rect 1029 -3439 1049 -1961
rect -1049 -3480 1049 -3439
rect 1449 -1961 3547 -1920
rect 1449 -3439 3291 -1961
rect 3527 -3439 3547 -1961
rect 1449 -3480 3547 -3439
rect 3947 -1961 6045 -1920
rect 3947 -3439 5789 -1961
rect 6025 -3439 6045 -1961
rect 3947 -3480 6045 -3439
rect 6445 -1961 8543 -1920
rect 6445 -3439 8287 -1961
rect 8523 -3439 8543 -1961
rect 6445 -3480 8543 -3439
rect 8943 -1961 11041 -1920
rect 8943 -3439 10785 -1961
rect 11021 -3439 11041 -1961
rect 8943 -3480 11041 -3439
rect -11041 -3761 -8943 -3720
rect -11041 -5239 -9199 -3761
rect -8963 -5239 -8943 -3761
rect -11041 -5280 -8943 -5239
rect -8543 -3761 -6445 -3720
rect -8543 -5239 -6701 -3761
rect -6465 -5239 -6445 -3761
rect -8543 -5280 -6445 -5239
rect -6045 -3761 -3947 -3720
rect -6045 -5239 -4203 -3761
rect -3967 -5239 -3947 -3761
rect -6045 -5280 -3947 -5239
rect -3547 -3761 -1449 -3720
rect -3547 -5239 -1705 -3761
rect -1469 -5239 -1449 -3761
rect -3547 -5280 -1449 -5239
rect -1049 -3761 1049 -3720
rect -1049 -5239 793 -3761
rect 1029 -5239 1049 -3761
rect -1049 -5280 1049 -5239
rect 1449 -3761 3547 -3720
rect 1449 -5239 3291 -3761
rect 3527 -5239 3547 -3761
rect 1449 -5280 3547 -5239
rect 3947 -3761 6045 -3720
rect 3947 -5239 5789 -3761
rect 6025 -5239 6045 -3761
rect 3947 -5280 6045 -5239
rect 6445 -3761 8543 -3720
rect 6445 -5239 8287 -3761
rect 8523 -5239 8543 -3761
rect 6445 -5280 8543 -5239
rect 8943 -3761 11041 -3720
rect 8943 -5239 10785 -3761
rect 11021 -5239 11041 -3761
rect 8943 -5280 11041 -5239
rect -11041 -5561 -8943 -5520
rect -11041 -7039 -9199 -5561
rect -8963 -7039 -8943 -5561
rect -11041 -7080 -8943 -7039
rect -8543 -5561 -6445 -5520
rect -8543 -7039 -6701 -5561
rect -6465 -7039 -6445 -5561
rect -8543 -7080 -6445 -7039
rect -6045 -5561 -3947 -5520
rect -6045 -7039 -4203 -5561
rect -3967 -7039 -3947 -5561
rect -6045 -7080 -3947 -7039
rect -3547 -5561 -1449 -5520
rect -3547 -7039 -1705 -5561
rect -1469 -7039 -1449 -5561
rect -3547 -7080 -1449 -7039
rect -1049 -5561 1049 -5520
rect -1049 -7039 793 -5561
rect 1029 -7039 1049 -5561
rect -1049 -7080 1049 -7039
rect 1449 -5561 3547 -5520
rect 1449 -7039 3291 -5561
rect 3527 -7039 3547 -5561
rect 1449 -7080 3547 -7039
rect 3947 -5561 6045 -5520
rect 3947 -7039 5789 -5561
rect 6025 -7039 6045 -5561
rect 3947 -7080 6045 -7039
rect 6445 -5561 8543 -5520
rect 6445 -7039 8287 -5561
rect 8523 -7039 8543 -5561
rect 6445 -7080 8543 -7039
rect 8943 -5561 11041 -5520
rect 8943 -7039 10785 -5561
rect 11021 -7039 11041 -5561
rect 8943 -7080 11041 -7039
rect -11041 -7361 -8943 -7320
rect -11041 -8839 -9199 -7361
rect -8963 -8839 -8943 -7361
rect -11041 -8880 -8943 -8839
rect -8543 -7361 -6445 -7320
rect -8543 -8839 -6701 -7361
rect -6465 -8839 -6445 -7361
rect -8543 -8880 -6445 -8839
rect -6045 -7361 -3947 -7320
rect -6045 -8839 -4203 -7361
rect -3967 -8839 -3947 -7361
rect -6045 -8880 -3947 -8839
rect -3547 -7361 -1449 -7320
rect -3547 -8839 -1705 -7361
rect -1469 -8839 -1449 -7361
rect -3547 -8880 -1449 -8839
rect -1049 -7361 1049 -7320
rect -1049 -8839 793 -7361
rect 1029 -8839 1049 -7361
rect -1049 -8880 1049 -8839
rect 1449 -7361 3547 -7320
rect 1449 -8839 3291 -7361
rect 3527 -8839 3547 -7361
rect 1449 -8880 3547 -8839
rect 3947 -7361 6045 -7320
rect 3947 -8839 5789 -7361
rect 6025 -8839 6045 -7361
rect 3947 -8880 6045 -8839
rect 6445 -7361 8543 -7320
rect 6445 -8839 8287 -7361
rect 8523 -8839 8543 -7361
rect 6445 -8880 8543 -8839
rect 8943 -7361 11041 -7320
rect 8943 -8839 10785 -7361
rect 11021 -8839 11041 -7361
rect 8943 -8880 11041 -8839
<< via4 >>
rect -9199 7361 -8963 8839
rect -6701 7361 -6465 8839
rect -4203 7361 -3967 8839
rect -1705 7361 -1469 8839
rect 793 7361 1029 8839
rect 3291 7361 3527 8839
rect 5789 7361 6025 8839
rect 8287 7361 8523 8839
rect 10785 7361 11021 8839
rect -9199 5561 -8963 7039
rect -6701 5561 -6465 7039
rect -4203 5561 -3967 7039
rect -1705 5561 -1469 7039
rect 793 5561 1029 7039
rect 3291 5561 3527 7039
rect 5789 5561 6025 7039
rect 8287 5561 8523 7039
rect 10785 5561 11021 7039
rect -9199 3761 -8963 5239
rect -6701 3761 -6465 5239
rect -4203 3761 -3967 5239
rect -1705 3761 -1469 5239
rect 793 3761 1029 5239
rect 3291 3761 3527 5239
rect 5789 3761 6025 5239
rect 8287 3761 8523 5239
rect 10785 3761 11021 5239
rect -9199 1961 -8963 3439
rect -6701 1961 -6465 3439
rect -4203 1961 -3967 3439
rect -1705 1961 -1469 3439
rect 793 1961 1029 3439
rect 3291 1961 3527 3439
rect 5789 1961 6025 3439
rect 8287 1961 8523 3439
rect 10785 1961 11021 3439
rect -9199 161 -8963 1639
rect -6701 161 -6465 1639
rect -4203 161 -3967 1639
rect -1705 161 -1469 1639
rect 793 161 1029 1639
rect 3291 161 3527 1639
rect 5789 161 6025 1639
rect 8287 161 8523 1639
rect 10785 161 11021 1639
rect -9199 -1639 -8963 -161
rect -6701 -1639 -6465 -161
rect -4203 -1639 -3967 -161
rect -1705 -1639 -1469 -161
rect 793 -1639 1029 -161
rect 3291 -1639 3527 -161
rect 5789 -1639 6025 -161
rect 8287 -1639 8523 -161
rect 10785 -1639 11021 -161
rect -9199 -3439 -8963 -1961
rect -6701 -3439 -6465 -1961
rect -4203 -3439 -3967 -1961
rect -1705 -3439 -1469 -1961
rect 793 -3439 1029 -1961
rect 3291 -3439 3527 -1961
rect 5789 -3439 6025 -1961
rect 8287 -3439 8523 -1961
rect 10785 -3439 11021 -1961
rect -9199 -5239 -8963 -3761
rect -6701 -5239 -6465 -3761
rect -4203 -5239 -3967 -3761
rect -1705 -5239 -1469 -3761
rect 793 -5239 1029 -3761
rect 3291 -5239 3527 -3761
rect 5789 -5239 6025 -3761
rect 8287 -5239 8523 -3761
rect 10785 -5239 11021 -3761
rect -9199 -7039 -8963 -5561
rect -6701 -7039 -6465 -5561
rect -4203 -7039 -3967 -5561
rect -1705 -7039 -1469 -5561
rect 793 -7039 1029 -5561
rect 3291 -7039 3527 -5561
rect 5789 -7039 6025 -5561
rect 8287 -7039 8523 -5561
rect 10785 -7039 11021 -5561
rect -9199 -8839 -8963 -7361
rect -6701 -8839 -6465 -7361
rect -4203 -8839 -3967 -7361
rect -1705 -8839 -1469 -7361
rect 793 -8839 1029 -7361
rect 3291 -8839 3527 -7361
rect 5789 -8839 6025 -7361
rect 8287 -8839 8523 -7361
rect 10785 -8839 11021 -7361
<< mimcap2 >>
rect -10961 8760 -9561 8800
rect -10961 7440 -10921 8760
rect -9601 7440 -9561 8760
rect -10961 7400 -9561 7440
rect -8463 8760 -7063 8800
rect -8463 7440 -8423 8760
rect -7103 7440 -7063 8760
rect -8463 7400 -7063 7440
rect -5965 8760 -4565 8800
rect -5965 7440 -5925 8760
rect -4605 7440 -4565 8760
rect -5965 7400 -4565 7440
rect -3467 8760 -2067 8800
rect -3467 7440 -3427 8760
rect -2107 7440 -2067 8760
rect -3467 7400 -2067 7440
rect -969 8760 431 8800
rect -969 7440 -929 8760
rect 391 7440 431 8760
rect -969 7400 431 7440
rect 1529 8760 2929 8800
rect 1529 7440 1569 8760
rect 2889 7440 2929 8760
rect 1529 7400 2929 7440
rect 4027 8760 5427 8800
rect 4027 7440 4067 8760
rect 5387 7440 5427 8760
rect 4027 7400 5427 7440
rect 6525 8760 7925 8800
rect 6525 7440 6565 8760
rect 7885 7440 7925 8760
rect 6525 7400 7925 7440
rect 9023 8760 10423 8800
rect 9023 7440 9063 8760
rect 10383 7440 10423 8760
rect 9023 7400 10423 7440
rect -10961 6960 -9561 7000
rect -10961 5640 -10921 6960
rect -9601 5640 -9561 6960
rect -10961 5600 -9561 5640
rect -8463 6960 -7063 7000
rect -8463 5640 -8423 6960
rect -7103 5640 -7063 6960
rect -8463 5600 -7063 5640
rect -5965 6960 -4565 7000
rect -5965 5640 -5925 6960
rect -4605 5640 -4565 6960
rect -5965 5600 -4565 5640
rect -3467 6960 -2067 7000
rect -3467 5640 -3427 6960
rect -2107 5640 -2067 6960
rect -3467 5600 -2067 5640
rect -969 6960 431 7000
rect -969 5640 -929 6960
rect 391 5640 431 6960
rect -969 5600 431 5640
rect 1529 6960 2929 7000
rect 1529 5640 1569 6960
rect 2889 5640 2929 6960
rect 1529 5600 2929 5640
rect 4027 6960 5427 7000
rect 4027 5640 4067 6960
rect 5387 5640 5427 6960
rect 4027 5600 5427 5640
rect 6525 6960 7925 7000
rect 6525 5640 6565 6960
rect 7885 5640 7925 6960
rect 6525 5600 7925 5640
rect 9023 6960 10423 7000
rect 9023 5640 9063 6960
rect 10383 5640 10423 6960
rect 9023 5600 10423 5640
rect -10961 5160 -9561 5200
rect -10961 3840 -10921 5160
rect -9601 3840 -9561 5160
rect -10961 3800 -9561 3840
rect -8463 5160 -7063 5200
rect -8463 3840 -8423 5160
rect -7103 3840 -7063 5160
rect -8463 3800 -7063 3840
rect -5965 5160 -4565 5200
rect -5965 3840 -5925 5160
rect -4605 3840 -4565 5160
rect -5965 3800 -4565 3840
rect -3467 5160 -2067 5200
rect -3467 3840 -3427 5160
rect -2107 3840 -2067 5160
rect -3467 3800 -2067 3840
rect -969 5160 431 5200
rect -969 3840 -929 5160
rect 391 3840 431 5160
rect -969 3800 431 3840
rect 1529 5160 2929 5200
rect 1529 3840 1569 5160
rect 2889 3840 2929 5160
rect 1529 3800 2929 3840
rect 4027 5160 5427 5200
rect 4027 3840 4067 5160
rect 5387 3840 5427 5160
rect 4027 3800 5427 3840
rect 6525 5160 7925 5200
rect 6525 3840 6565 5160
rect 7885 3840 7925 5160
rect 6525 3800 7925 3840
rect 9023 5160 10423 5200
rect 9023 3840 9063 5160
rect 10383 3840 10423 5160
rect 9023 3800 10423 3840
rect -10961 3360 -9561 3400
rect -10961 2040 -10921 3360
rect -9601 2040 -9561 3360
rect -10961 2000 -9561 2040
rect -8463 3360 -7063 3400
rect -8463 2040 -8423 3360
rect -7103 2040 -7063 3360
rect -8463 2000 -7063 2040
rect -5965 3360 -4565 3400
rect -5965 2040 -5925 3360
rect -4605 2040 -4565 3360
rect -5965 2000 -4565 2040
rect -3467 3360 -2067 3400
rect -3467 2040 -3427 3360
rect -2107 2040 -2067 3360
rect -3467 2000 -2067 2040
rect -969 3360 431 3400
rect -969 2040 -929 3360
rect 391 2040 431 3360
rect -969 2000 431 2040
rect 1529 3360 2929 3400
rect 1529 2040 1569 3360
rect 2889 2040 2929 3360
rect 1529 2000 2929 2040
rect 4027 3360 5427 3400
rect 4027 2040 4067 3360
rect 5387 2040 5427 3360
rect 4027 2000 5427 2040
rect 6525 3360 7925 3400
rect 6525 2040 6565 3360
rect 7885 2040 7925 3360
rect 6525 2000 7925 2040
rect 9023 3360 10423 3400
rect 9023 2040 9063 3360
rect 10383 2040 10423 3360
rect 9023 2000 10423 2040
rect -10961 1560 -9561 1600
rect -10961 240 -10921 1560
rect -9601 240 -9561 1560
rect -10961 200 -9561 240
rect -8463 1560 -7063 1600
rect -8463 240 -8423 1560
rect -7103 240 -7063 1560
rect -8463 200 -7063 240
rect -5965 1560 -4565 1600
rect -5965 240 -5925 1560
rect -4605 240 -4565 1560
rect -5965 200 -4565 240
rect -3467 1560 -2067 1600
rect -3467 240 -3427 1560
rect -2107 240 -2067 1560
rect -3467 200 -2067 240
rect -969 1560 431 1600
rect -969 240 -929 1560
rect 391 240 431 1560
rect -969 200 431 240
rect 1529 1560 2929 1600
rect 1529 240 1569 1560
rect 2889 240 2929 1560
rect 1529 200 2929 240
rect 4027 1560 5427 1600
rect 4027 240 4067 1560
rect 5387 240 5427 1560
rect 4027 200 5427 240
rect 6525 1560 7925 1600
rect 6525 240 6565 1560
rect 7885 240 7925 1560
rect 6525 200 7925 240
rect 9023 1560 10423 1600
rect 9023 240 9063 1560
rect 10383 240 10423 1560
rect 9023 200 10423 240
rect -10961 -240 -9561 -200
rect -10961 -1560 -10921 -240
rect -9601 -1560 -9561 -240
rect -10961 -1600 -9561 -1560
rect -8463 -240 -7063 -200
rect -8463 -1560 -8423 -240
rect -7103 -1560 -7063 -240
rect -8463 -1600 -7063 -1560
rect -5965 -240 -4565 -200
rect -5965 -1560 -5925 -240
rect -4605 -1560 -4565 -240
rect -5965 -1600 -4565 -1560
rect -3467 -240 -2067 -200
rect -3467 -1560 -3427 -240
rect -2107 -1560 -2067 -240
rect -3467 -1600 -2067 -1560
rect -969 -240 431 -200
rect -969 -1560 -929 -240
rect 391 -1560 431 -240
rect -969 -1600 431 -1560
rect 1529 -240 2929 -200
rect 1529 -1560 1569 -240
rect 2889 -1560 2929 -240
rect 1529 -1600 2929 -1560
rect 4027 -240 5427 -200
rect 4027 -1560 4067 -240
rect 5387 -1560 5427 -240
rect 4027 -1600 5427 -1560
rect 6525 -240 7925 -200
rect 6525 -1560 6565 -240
rect 7885 -1560 7925 -240
rect 6525 -1600 7925 -1560
rect 9023 -240 10423 -200
rect 9023 -1560 9063 -240
rect 10383 -1560 10423 -240
rect 9023 -1600 10423 -1560
rect -10961 -2040 -9561 -2000
rect -10961 -3360 -10921 -2040
rect -9601 -3360 -9561 -2040
rect -10961 -3400 -9561 -3360
rect -8463 -2040 -7063 -2000
rect -8463 -3360 -8423 -2040
rect -7103 -3360 -7063 -2040
rect -8463 -3400 -7063 -3360
rect -5965 -2040 -4565 -2000
rect -5965 -3360 -5925 -2040
rect -4605 -3360 -4565 -2040
rect -5965 -3400 -4565 -3360
rect -3467 -2040 -2067 -2000
rect -3467 -3360 -3427 -2040
rect -2107 -3360 -2067 -2040
rect -3467 -3400 -2067 -3360
rect -969 -2040 431 -2000
rect -969 -3360 -929 -2040
rect 391 -3360 431 -2040
rect -969 -3400 431 -3360
rect 1529 -2040 2929 -2000
rect 1529 -3360 1569 -2040
rect 2889 -3360 2929 -2040
rect 1529 -3400 2929 -3360
rect 4027 -2040 5427 -2000
rect 4027 -3360 4067 -2040
rect 5387 -3360 5427 -2040
rect 4027 -3400 5427 -3360
rect 6525 -2040 7925 -2000
rect 6525 -3360 6565 -2040
rect 7885 -3360 7925 -2040
rect 6525 -3400 7925 -3360
rect 9023 -2040 10423 -2000
rect 9023 -3360 9063 -2040
rect 10383 -3360 10423 -2040
rect 9023 -3400 10423 -3360
rect -10961 -3840 -9561 -3800
rect -10961 -5160 -10921 -3840
rect -9601 -5160 -9561 -3840
rect -10961 -5200 -9561 -5160
rect -8463 -3840 -7063 -3800
rect -8463 -5160 -8423 -3840
rect -7103 -5160 -7063 -3840
rect -8463 -5200 -7063 -5160
rect -5965 -3840 -4565 -3800
rect -5965 -5160 -5925 -3840
rect -4605 -5160 -4565 -3840
rect -5965 -5200 -4565 -5160
rect -3467 -3840 -2067 -3800
rect -3467 -5160 -3427 -3840
rect -2107 -5160 -2067 -3840
rect -3467 -5200 -2067 -5160
rect -969 -3840 431 -3800
rect -969 -5160 -929 -3840
rect 391 -5160 431 -3840
rect -969 -5200 431 -5160
rect 1529 -3840 2929 -3800
rect 1529 -5160 1569 -3840
rect 2889 -5160 2929 -3840
rect 1529 -5200 2929 -5160
rect 4027 -3840 5427 -3800
rect 4027 -5160 4067 -3840
rect 5387 -5160 5427 -3840
rect 4027 -5200 5427 -5160
rect 6525 -3840 7925 -3800
rect 6525 -5160 6565 -3840
rect 7885 -5160 7925 -3840
rect 6525 -5200 7925 -5160
rect 9023 -3840 10423 -3800
rect 9023 -5160 9063 -3840
rect 10383 -5160 10423 -3840
rect 9023 -5200 10423 -5160
rect -10961 -5640 -9561 -5600
rect -10961 -6960 -10921 -5640
rect -9601 -6960 -9561 -5640
rect -10961 -7000 -9561 -6960
rect -8463 -5640 -7063 -5600
rect -8463 -6960 -8423 -5640
rect -7103 -6960 -7063 -5640
rect -8463 -7000 -7063 -6960
rect -5965 -5640 -4565 -5600
rect -5965 -6960 -5925 -5640
rect -4605 -6960 -4565 -5640
rect -5965 -7000 -4565 -6960
rect -3467 -5640 -2067 -5600
rect -3467 -6960 -3427 -5640
rect -2107 -6960 -2067 -5640
rect -3467 -7000 -2067 -6960
rect -969 -5640 431 -5600
rect -969 -6960 -929 -5640
rect 391 -6960 431 -5640
rect -969 -7000 431 -6960
rect 1529 -5640 2929 -5600
rect 1529 -6960 1569 -5640
rect 2889 -6960 2929 -5640
rect 1529 -7000 2929 -6960
rect 4027 -5640 5427 -5600
rect 4027 -6960 4067 -5640
rect 5387 -6960 5427 -5640
rect 4027 -7000 5427 -6960
rect 6525 -5640 7925 -5600
rect 6525 -6960 6565 -5640
rect 7885 -6960 7925 -5640
rect 6525 -7000 7925 -6960
rect 9023 -5640 10423 -5600
rect 9023 -6960 9063 -5640
rect 10383 -6960 10423 -5640
rect 9023 -7000 10423 -6960
rect -10961 -7440 -9561 -7400
rect -10961 -8760 -10921 -7440
rect -9601 -8760 -9561 -7440
rect -10961 -8800 -9561 -8760
rect -8463 -7440 -7063 -7400
rect -8463 -8760 -8423 -7440
rect -7103 -8760 -7063 -7440
rect -8463 -8800 -7063 -8760
rect -5965 -7440 -4565 -7400
rect -5965 -8760 -5925 -7440
rect -4605 -8760 -4565 -7440
rect -5965 -8800 -4565 -8760
rect -3467 -7440 -2067 -7400
rect -3467 -8760 -3427 -7440
rect -2107 -8760 -2067 -7440
rect -3467 -8800 -2067 -8760
rect -969 -7440 431 -7400
rect -969 -8760 -929 -7440
rect 391 -8760 431 -7440
rect -969 -8800 431 -8760
rect 1529 -7440 2929 -7400
rect 1529 -8760 1569 -7440
rect 2889 -8760 2929 -7440
rect 1529 -8800 2929 -8760
rect 4027 -7440 5427 -7400
rect 4027 -8760 4067 -7440
rect 5387 -8760 5427 -7440
rect 4027 -8800 5427 -8760
rect 6525 -7440 7925 -7400
rect 6525 -8760 6565 -7440
rect 7885 -8760 7925 -7440
rect 6525 -8800 7925 -8760
rect 9023 -7440 10423 -7400
rect 9023 -8760 9063 -7440
rect 10383 -8760 10423 -7440
rect 9023 -8800 10423 -8760
<< mimcap2contact >>
rect -10921 7440 -9601 8760
rect -8423 7440 -7103 8760
rect -5925 7440 -4605 8760
rect -3427 7440 -2107 8760
rect -929 7440 391 8760
rect 1569 7440 2889 8760
rect 4067 7440 5387 8760
rect 6565 7440 7885 8760
rect 9063 7440 10383 8760
rect -10921 5640 -9601 6960
rect -8423 5640 -7103 6960
rect -5925 5640 -4605 6960
rect -3427 5640 -2107 6960
rect -929 5640 391 6960
rect 1569 5640 2889 6960
rect 4067 5640 5387 6960
rect 6565 5640 7885 6960
rect 9063 5640 10383 6960
rect -10921 3840 -9601 5160
rect -8423 3840 -7103 5160
rect -5925 3840 -4605 5160
rect -3427 3840 -2107 5160
rect -929 3840 391 5160
rect 1569 3840 2889 5160
rect 4067 3840 5387 5160
rect 6565 3840 7885 5160
rect 9063 3840 10383 5160
rect -10921 2040 -9601 3360
rect -8423 2040 -7103 3360
rect -5925 2040 -4605 3360
rect -3427 2040 -2107 3360
rect -929 2040 391 3360
rect 1569 2040 2889 3360
rect 4067 2040 5387 3360
rect 6565 2040 7885 3360
rect 9063 2040 10383 3360
rect -10921 240 -9601 1560
rect -8423 240 -7103 1560
rect -5925 240 -4605 1560
rect -3427 240 -2107 1560
rect -929 240 391 1560
rect 1569 240 2889 1560
rect 4067 240 5387 1560
rect 6565 240 7885 1560
rect 9063 240 10383 1560
rect -10921 -1560 -9601 -240
rect -8423 -1560 -7103 -240
rect -5925 -1560 -4605 -240
rect -3427 -1560 -2107 -240
rect -929 -1560 391 -240
rect 1569 -1560 2889 -240
rect 4067 -1560 5387 -240
rect 6565 -1560 7885 -240
rect 9063 -1560 10383 -240
rect -10921 -3360 -9601 -2040
rect -8423 -3360 -7103 -2040
rect -5925 -3360 -4605 -2040
rect -3427 -3360 -2107 -2040
rect -929 -3360 391 -2040
rect 1569 -3360 2889 -2040
rect 4067 -3360 5387 -2040
rect 6565 -3360 7885 -2040
rect 9063 -3360 10383 -2040
rect -10921 -5160 -9601 -3840
rect -8423 -5160 -7103 -3840
rect -5925 -5160 -4605 -3840
rect -3427 -5160 -2107 -3840
rect -929 -5160 391 -3840
rect 1569 -5160 2889 -3840
rect 4067 -5160 5387 -3840
rect 6565 -5160 7885 -3840
rect 9063 -5160 10383 -3840
rect -10921 -6960 -9601 -5640
rect -8423 -6960 -7103 -5640
rect -5925 -6960 -4605 -5640
rect -3427 -6960 -2107 -5640
rect -929 -6960 391 -5640
rect 1569 -6960 2889 -5640
rect 4067 -6960 5387 -5640
rect 6565 -6960 7885 -5640
rect 9063 -6960 10383 -5640
rect -10921 -8760 -9601 -7440
rect -8423 -8760 -7103 -7440
rect -5925 -8760 -4605 -7440
rect -3427 -8760 -2107 -7440
rect -929 -8760 391 -7440
rect 1569 -8760 2889 -7440
rect 4067 -8760 5387 -7440
rect 6565 -8760 7885 -7440
rect 9063 -8760 10383 -7440
<< metal5 >>
rect -9241 8839 -8921 8881
rect -10945 8760 -9577 8784
rect -10945 7440 -10921 8760
rect -9601 7440 -9577 8760
rect -10945 7416 -9577 7440
rect -9241 7361 -9199 8839
rect -8963 7361 -8921 8839
rect -6743 8839 -6423 8881
rect -8447 8760 -7079 8784
rect -8447 7440 -8423 8760
rect -7103 7440 -7079 8760
rect -8447 7416 -7079 7440
rect -9241 7319 -8921 7361
rect -6743 7361 -6701 8839
rect -6465 7361 -6423 8839
rect -4245 8839 -3925 8881
rect -5949 8760 -4581 8784
rect -5949 7440 -5925 8760
rect -4605 7440 -4581 8760
rect -5949 7416 -4581 7440
rect -6743 7319 -6423 7361
rect -4245 7361 -4203 8839
rect -3967 7361 -3925 8839
rect -1747 8839 -1427 8881
rect -3451 8760 -2083 8784
rect -3451 7440 -3427 8760
rect -2107 7440 -2083 8760
rect -3451 7416 -2083 7440
rect -4245 7319 -3925 7361
rect -1747 7361 -1705 8839
rect -1469 7361 -1427 8839
rect 751 8839 1071 8881
rect -953 8760 415 8784
rect -953 7440 -929 8760
rect 391 7440 415 8760
rect -953 7416 415 7440
rect -1747 7319 -1427 7361
rect 751 7361 793 8839
rect 1029 7361 1071 8839
rect 3249 8839 3569 8881
rect 1545 8760 2913 8784
rect 1545 7440 1569 8760
rect 2889 7440 2913 8760
rect 1545 7416 2913 7440
rect 751 7319 1071 7361
rect 3249 7361 3291 8839
rect 3527 7361 3569 8839
rect 5747 8839 6067 8881
rect 4043 8760 5411 8784
rect 4043 7440 4067 8760
rect 5387 7440 5411 8760
rect 4043 7416 5411 7440
rect 3249 7319 3569 7361
rect 5747 7361 5789 8839
rect 6025 7361 6067 8839
rect 8245 8839 8565 8881
rect 6541 8760 7909 8784
rect 6541 7440 6565 8760
rect 7885 7440 7909 8760
rect 6541 7416 7909 7440
rect 5747 7319 6067 7361
rect 8245 7361 8287 8839
rect 8523 7361 8565 8839
rect 10743 8839 11063 8881
rect 9039 8760 10407 8784
rect 9039 7440 9063 8760
rect 10383 7440 10407 8760
rect 9039 7416 10407 7440
rect 8245 7319 8565 7361
rect 10743 7361 10785 8839
rect 11021 7361 11063 8839
rect 10743 7319 11063 7361
rect -9241 7039 -8921 7081
rect -10945 6960 -9577 6984
rect -10945 5640 -10921 6960
rect -9601 5640 -9577 6960
rect -10945 5616 -9577 5640
rect -9241 5561 -9199 7039
rect -8963 5561 -8921 7039
rect -6743 7039 -6423 7081
rect -8447 6960 -7079 6984
rect -8447 5640 -8423 6960
rect -7103 5640 -7079 6960
rect -8447 5616 -7079 5640
rect -9241 5519 -8921 5561
rect -6743 5561 -6701 7039
rect -6465 5561 -6423 7039
rect -4245 7039 -3925 7081
rect -5949 6960 -4581 6984
rect -5949 5640 -5925 6960
rect -4605 5640 -4581 6960
rect -5949 5616 -4581 5640
rect -6743 5519 -6423 5561
rect -4245 5561 -4203 7039
rect -3967 5561 -3925 7039
rect -1747 7039 -1427 7081
rect -3451 6960 -2083 6984
rect -3451 5640 -3427 6960
rect -2107 5640 -2083 6960
rect -3451 5616 -2083 5640
rect -4245 5519 -3925 5561
rect -1747 5561 -1705 7039
rect -1469 5561 -1427 7039
rect 751 7039 1071 7081
rect -953 6960 415 6984
rect -953 5640 -929 6960
rect 391 5640 415 6960
rect -953 5616 415 5640
rect -1747 5519 -1427 5561
rect 751 5561 793 7039
rect 1029 5561 1071 7039
rect 3249 7039 3569 7081
rect 1545 6960 2913 6984
rect 1545 5640 1569 6960
rect 2889 5640 2913 6960
rect 1545 5616 2913 5640
rect 751 5519 1071 5561
rect 3249 5561 3291 7039
rect 3527 5561 3569 7039
rect 5747 7039 6067 7081
rect 4043 6960 5411 6984
rect 4043 5640 4067 6960
rect 5387 5640 5411 6960
rect 4043 5616 5411 5640
rect 3249 5519 3569 5561
rect 5747 5561 5789 7039
rect 6025 5561 6067 7039
rect 8245 7039 8565 7081
rect 6541 6960 7909 6984
rect 6541 5640 6565 6960
rect 7885 5640 7909 6960
rect 6541 5616 7909 5640
rect 5747 5519 6067 5561
rect 8245 5561 8287 7039
rect 8523 5561 8565 7039
rect 10743 7039 11063 7081
rect 9039 6960 10407 6984
rect 9039 5640 9063 6960
rect 10383 5640 10407 6960
rect 9039 5616 10407 5640
rect 8245 5519 8565 5561
rect 10743 5561 10785 7039
rect 11021 5561 11063 7039
rect 10743 5519 11063 5561
rect -9241 5239 -8921 5281
rect -10945 5160 -9577 5184
rect -10945 3840 -10921 5160
rect -9601 3840 -9577 5160
rect -10945 3816 -9577 3840
rect -9241 3761 -9199 5239
rect -8963 3761 -8921 5239
rect -6743 5239 -6423 5281
rect -8447 5160 -7079 5184
rect -8447 3840 -8423 5160
rect -7103 3840 -7079 5160
rect -8447 3816 -7079 3840
rect -9241 3719 -8921 3761
rect -6743 3761 -6701 5239
rect -6465 3761 -6423 5239
rect -4245 5239 -3925 5281
rect -5949 5160 -4581 5184
rect -5949 3840 -5925 5160
rect -4605 3840 -4581 5160
rect -5949 3816 -4581 3840
rect -6743 3719 -6423 3761
rect -4245 3761 -4203 5239
rect -3967 3761 -3925 5239
rect -1747 5239 -1427 5281
rect -3451 5160 -2083 5184
rect -3451 3840 -3427 5160
rect -2107 3840 -2083 5160
rect -3451 3816 -2083 3840
rect -4245 3719 -3925 3761
rect -1747 3761 -1705 5239
rect -1469 3761 -1427 5239
rect 751 5239 1071 5281
rect -953 5160 415 5184
rect -953 3840 -929 5160
rect 391 3840 415 5160
rect -953 3816 415 3840
rect -1747 3719 -1427 3761
rect 751 3761 793 5239
rect 1029 3761 1071 5239
rect 3249 5239 3569 5281
rect 1545 5160 2913 5184
rect 1545 3840 1569 5160
rect 2889 3840 2913 5160
rect 1545 3816 2913 3840
rect 751 3719 1071 3761
rect 3249 3761 3291 5239
rect 3527 3761 3569 5239
rect 5747 5239 6067 5281
rect 4043 5160 5411 5184
rect 4043 3840 4067 5160
rect 5387 3840 5411 5160
rect 4043 3816 5411 3840
rect 3249 3719 3569 3761
rect 5747 3761 5789 5239
rect 6025 3761 6067 5239
rect 8245 5239 8565 5281
rect 6541 5160 7909 5184
rect 6541 3840 6565 5160
rect 7885 3840 7909 5160
rect 6541 3816 7909 3840
rect 5747 3719 6067 3761
rect 8245 3761 8287 5239
rect 8523 3761 8565 5239
rect 10743 5239 11063 5281
rect 9039 5160 10407 5184
rect 9039 3840 9063 5160
rect 10383 3840 10407 5160
rect 9039 3816 10407 3840
rect 8245 3719 8565 3761
rect 10743 3761 10785 5239
rect 11021 3761 11063 5239
rect 10743 3719 11063 3761
rect -9241 3439 -8921 3481
rect -10945 3360 -9577 3384
rect -10945 2040 -10921 3360
rect -9601 2040 -9577 3360
rect -10945 2016 -9577 2040
rect -9241 1961 -9199 3439
rect -8963 1961 -8921 3439
rect -6743 3439 -6423 3481
rect -8447 3360 -7079 3384
rect -8447 2040 -8423 3360
rect -7103 2040 -7079 3360
rect -8447 2016 -7079 2040
rect -9241 1919 -8921 1961
rect -6743 1961 -6701 3439
rect -6465 1961 -6423 3439
rect -4245 3439 -3925 3481
rect -5949 3360 -4581 3384
rect -5949 2040 -5925 3360
rect -4605 2040 -4581 3360
rect -5949 2016 -4581 2040
rect -6743 1919 -6423 1961
rect -4245 1961 -4203 3439
rect -3967 1961 -3925 3439
rect -1747 3439 -1427 3481
rect -3451 3360 -2083 3384
rect -3451 2040 -3427 3360
rect -2107 2040 -2083 3360
rect -3451 2016 -2083 2040
rect -4245 1919 -3925 1961
rect -1747 1961 -1705 3439
rect -1469 1961 -1427 3439
rect 751 3439 1071 3481
rect -953 3360 415 3384
rect -953 2040 -929 3360
rect 391 2040 415 3360
rect -953 2016 415 2040
rect -1747 1919 -1427 1961
rect 751 1961 793 3439
rect 1029 1961 1071 3439
rect 3249 3439 3569 3481
rect 1545 3360 2913 3384
rect 1545 2040 1569 3360
rect 2889 2040 2913 3360
rect 1545 2016 2913 2040
rect 751 1919 1071 1961
rect 3249 1961 3291 3439
rect 3527 1961 3569 3439
rect 5747 3439 6067 3481
rect 4043 3360 5411 3384
rect 4043 2040 4067 3360
rect 5387 2040 5411 3360
rect 4043 2016 5411 2040
rect 3249 1919 3569 1961
rect 5747 1961 5789 3439
rect 6025 1961 6067 3439
rect 8245 3439 8565 3481
rect 6541 3360 7909 3384
rect 6541 2040 6565 3360
rect 7885 2040 7909 3360
rect 6541 2016 7909 2040
rect 5747 1919 6067 1961
rect 8245 1961 8287 3439
rect 8523 1961 8565 3439
rect 10743 3439 11063 3481
rect 9039 3360 10407 3384
rect 9039 2040 9063 3360
rect 10383 2040 10407 3360
rect 9039 2016 10407 2040
rect 8245 1919 8565 1961
rect 10743 1961 10785 3439
rect 11021 1961 11063 3439
rect 10743 1919 11063 1961
rect -9241 1639 -8921 1681
rect -10945 1560 -9577 1584
rect -10945 240 -10921 1560
rect -9601 240 -9577 1560
rect -10945 216 -9577 240
rect -9241 161 -9199 1639
rect -8963 161 -8921 1639
rect -6743 1639 -6423 1681
rect -8447 1560 -7079 1584
rect -8447 240 -8423 1560
rect -7103 240 -7079 1560
rect -8447 216 -7079 240
rect -9241 119 -8921 161
rect -6743 161 -6701 1639
rect -6465 161 -6423 1639
rect -4245 1639 -3925 1681
rect -5949 1560 -4581 1584
rect -5949 240 -5925 1560
rect -4605 240 -4581 1560
rect -5949 216 -4581 240
rect -6743 119 -6423 161
rect -4245 161 -4203 1639
rect -3967 161 -3925 1639
rect -1747 1639 -1427 1681
rect -3451 1560 -2083 1584
rect -3451 240 -3427 1560
rect -2107 240 -2083 1560
rect -3451 216 -2083 240
rect -4245 119 -3925 161
rect -1747 161 -1705 1639
rect -1469 161 -1427 1639
rect 751 1639 1071 1681
rect -953 1560 415 1584
rect -953 240 -929 1560
rect 391 240 415 1560
rect -953 216 415 240
rect -1747 119 -1427 161
rect 751 161 793 1639
rect 1029 161 1071 1639
rect 3249 1639 3569 1681
rect 1545 1560 2913 1584
rect 1545 240 1569 1560
rect 2889 240 2913 1560
rect 1545 216 2913 240
rect 751 119 1071 161
rect 3249 161 3291 1639
rect 3527 161 3569 1639
rect 5747 1639 6067 1681
rect 4043 1560 5411 1584
rect 4043 240 4067 1560
rect 5387 240 5411 1560
rect 4043 216 5411 240
rect 3249 119 3569 161
rect 5747 161 5789 1639
rect 6025 161 6067 1639
rect 8245 1639 8565 1681
rect 6541 1560 7909 1584
rect 6541 240 6565 1560
rect 7885 240 7909 1560
rect 6541 216 7909 240
rect 5747 119 6067 161
rect 8245 161 8287 1639
rect 8523 161 8565 1639
rect 10743 1639 11063 1681
rect 9039 1560 10407 1584
rect 9039 240 9063 1560
rect 10383 240 10407 1560
rect 9039 216 10407 240
rect 8245 119 8565 161
rect 10743 161 10785 1639
rect 11021 161 11063 1639
rect 10743 119 11063 161
rect -9241 -161 -8921 -119
rect -10945 -240 -9577 -216
rect -10945 -1560 -10921 -240
rect -9601 -1560 -9577 -240
rect -10945 -1584 -9577 -1560
rect -9241 -1639 -9199 -161
rect -8963 -1639 -8921 -161
rect -6743 -161 -6423 -119
rect -8447 -240 -7079 -216
rect -8447 -1560 -8423 -240
rect -7103 -1560 -7079 -240
rect -8447 -1584 -7079 -1560
rect -9241 -1681 -8921 -1639
rect -6743 -1639 -6701 -161
rect -6465 -1639 -6423 -161
rect -4245 -161 -3925 -119
rect -5949 -240 -4581 -216
rect -5949 -1560 -5925 -240
rect -4605 -1560 -4581 -240
rect -5949 -1584 -4581 -1560
rect -6743 -1681 -6423 -1639
rect -4245 -1639 -4203 -161
rect -3967 -1639 -3925 -161
rect -1747 -161 -1427 -119
rect -3451 -240 -2083 -216
rect -3451 -1560 -3427 -240
rect -2107 -1560 -2083 -240
rect -3451 -1584 -2083 -1560
rect -4245 -1681 -3925 -1639
rect -1747 -1639 -1705 -161
rect -1469 -1639 -1427 -161
rect 751 -161 1071 -119
rect -953 -240 415 -216
rect -953 -1560 -929 -240
rect 391 -1560 415 -240
rect -953 -1584 415 -1560
rect -1747 -1681 -1427 -1639
rect 751 -1639 793 -161
rect 1029 -1639 1071 -161
rect 3249 -161 3569 -119
rect 1545 -240 2913 -216
rect 1545 -1560 1569 -240
rect 2889 -1560 2913 -240
rect 1545 -1584 2913 -1560
rect 751 -1681 1071 -1639
rect 3249 -1639 3291 -161
rect 3527 -1639 3569 -161
rect 5747 -161 6067 -119
rect 4043 -240 5411 -216
rect 4043 -1560 4067 -240
rect 5387 -1560 5411 -240
rect 4043 -1584 5411 -1560
rect 3249 -1681 3569 -1639
rect 5747 -1639 5789 -161
rect 6025 -1639 6067 -161
rect 8245 -161 8565 -119
rect 6541 -240 7909 -216
rect 6541 -1560 6565 -240
rect 7885 -1560 7909 -240
rect 6541 -1584 7909 -1560
rect 5747 -1681 6067 -1639
rect 8245 -1639 8287 -161
rect 8523 -1639 8565 -161
rect 10743 -161 11063 -119
rect 9039 -240 10407 -216
rect 9039 -1560 9063 -240
rect 10383 -1560 10407 -240
rect 9039 -1584 10407 -1560
rect 8245 -1681 8565 -1639
rect 10743 -1639 10785 -161
rect 11021 -1639 11063 -161
rect 10743 -1681 11063 -1639
rect -9241 -1961 -8921 -1919
rect -10945 -2040 -9577 -2016
rect -10945 -3360 -10921 -2040
rect -9601 -3360 -9577 -2040
rect -10945 -3384 -9577 -3360
rect -9241 -3439 -9199 -1961
rect -8963 -3439 -8921 -1961
rect -6743 -1961 -6423 -1919
rect -8447 -2040 -7079 -2016
rect -8447 -3360 -8423 -2040
rect -7103 -3360 -7079 -2040
rect -8447 -3384 -7079 -3360
rect -9241 -3481 -8921 -3439
rect -6743 -3439 -6701 -1961
rect -6465 -3439 -6423 -1961
rect -4245 -1961 -3925 -1919
rect -5949 -2040 -4581 -2016
rect -5949 -3360 -5925 -2040
rect -4605 -3360 -4581 -2040
rect -5949 -3384 -4581 -3360
rect -6743 -3481 -6423 -3439
rect -4245 -3439 -4203 -1961
rect -3967 -3439 -3925 -1961
rect -1747 -1961 -1427 -1919
rect -3451 -2040 -2083 -2016
rect -3451 -3360 -3427 -2040
rect -2107 -3360 -2083 -2040
rect -3451 -3384 -2083 -3360
rect -4245 -3481 -3925 -3439
rect -1747 -3439 -1705 -1961
rect -1469 -3439 -1427 -1961
rect 751 -1961 1071 -1919
rect -953 -2040 415 -2016
rect -953 -3360 -929 -2040
rect 391 -3360 415 -2040
rect -953 -3384 415 -3360
rect -1747 -3481 -1427 -3439
rect 751 -3439 793 -1961
rect 1029 -3439 1071 -1961
rect 3249 -1961 3569 -1919
rect 1545 -2040 2913 -2016
rect 1545 -3360 1569 -2040
rect 2889 -3360 2913 -2040
rect 1545 -3384 2913 -3360
rect 751 -3481 1071 -3439
rect 3249 -3439 3291 -1961
rect 3527 -3439 3569 -1961
rect 5747 -1961 6067 -1919
rect 4043 -2040 5411 -2016
rect 4043 -3360 4067 -2040
rect 5387 -3360 5411 -2040
rect 4043 -3384 5411 -3360
rect 3249 -3481 3569 -3439
rect 5747 -3439 5789 -1961
rect 6025 -3439 6067 -1961
rect 8245 -1961 8565 -1919
rect 6541 -2040 7909 -2016
rect 6541 -3360 6565 -2040
rect 7885 -3360 7909 -2040
rect 6541 -3384 7909 -3360
rect 5747 -3481 6067 -3439
rect 8245 -3439 8287 -1961
rect 8523 -3439 8565 -1961
rect 10743 -1961 11063 -1919
rect 9039 -2040 10407 -2016
rect 9039 -3360 9063 -2040
rect 10383 -3360 10407 -2040
rect 9039 -3384 10407 -3360
rect 8245 -3481 8565 -3439
rect 10743 -3439 10785 -1961
rect 11021 -3439 11063 -1961
rect 10743 -3481 11063 -3439
rect -9241 -3761 -8921 -3719
rect -10945 -3840 -9577 -3816
rect -10945 -5160 -10921 -3840
rect -9601 -5160 -9577 -3840
rect -10945 -5184 -9577 -5160
rect -9241 -5239 -9199 -3761
rect -8963 -5239 -8921 -3761
rect -6743 -3761 -6423 -3719
rect -8447 -3840 -7079 -3816
rect -8447 -5160 -8423 -3840
rect -7103 -5160 -7079 -3840
rect -8447 -5184 -7079 -5160
rect -9241 -5281 -8921 -5239
rect -6743 -5239 -6701 -3761
rect -6465 -5239 -6423 -3761
rect -4245 -3761 -3925 -3719
rect -5949 -3840 -4581 -3816
rect -5949 -5160 -5925 -3840
rect -4605 -5160 -4581 -3840
rect -5949 -5184 -4581 -5160
rect -6743 -5281 -6423 -5239
rect -4245 -5239 -4203 -3761
rect -3967 -5239 -3925 -3761
rect -1747 -3761 -1427 -3719
rect -3451 -3840 -2083 -3816
rect -3451 -5160 -3427 -3840
rect -2107 -5160 -2083 -3840
rect -3451 -5184 -2083 -5160
rect -4245 -5281 -3925 -5239
rect -1747 -5239 -1705 -3761
rect -1469 -5239 -1427 -3761
rect 751 -3761 1071 -3719
rect -953 -3840 415 -3816
rect -953 -5160 -929 -3840
rect 391 -5160 415 -3840
rect -953 -5184 415 -5160
rect -1747 -5281 -1427 -5239
rect 751 -5239 793 -3761
rect 1029 -5239 1071 -3761
rect 3249 -3761 3569 -3719
rect 1545 -3840 2913 -3816
rect 1545 -5160 1569 -3840
rect 2889 -5160 2913 -3840
rect 1545 -5184 2913 -5160
rect 751 -5281 1071 -5239
rect 3249 -5239 3291 -3761
rect 3527 -5239 3569 -3761
rect 5747 -3761 6067 -3719
rect 4043 -3840 5411 -3816
rect 4043 -5160 4067 -3840
rect 5387 -5160 5411 -3840
rect 4043 -5184 5411 -5160
rect 3249 -5281 3569 -5239
rect 5747 -5239 5789 -3761
rect 6025 -5239 6067 -3761
rect 8245 -3761 8565 -3719
rect 6541 -3840 7909 -3816
rect 6541 -5160 6565 -3840
rect 7885 -5160 7909 -3840
rect 6541 -5184 7909 -5160
rect 5747 -5281 6067 -5239
rect 8245 -5239 8287 -3761
rect 8523 -5239 8565 -3761
rect 10743 -3761 11063 -3719
rect 9039 -3840 10407 -3816
rect 9039 -5160 9063 -3840
rect 10383 -5160 10407 -3840
rect 9039 -5184 10407 -5160
rect 8245 -5281 8565 -5239
rect 10743 -5239 10785 -3761
rect 11021 -5239 11063 -3761
rect 10743 -5281 11063 -5239
rect -9241 -5561 -8921 -5519
rect -10945 -5640 -9577 -5616
rect -10945 -6960 -10921 -5640
rect -9601 -6960 -9577 -5640
rect -10945 -6984 -9577 -6960
rect -9241 -7039 -9199 -5561
rect -8963 -7039 -8921 -5561
rect -6743 -5561 -6423 -5519
rect -8447 -5640 -7079 -5616
rect -8447 -6960 -8423 -5640
rect -7103 -6960 -7079 -5640
rect -8447 -6984 -7079 -6960
rect -9241 -7081 -8921 -7039
rect -6743 -7039 -6701 -5561
rect -6465 -7039 -6423 -5561
rect -4245 -5561 -3925 -5519
rect -5949 -5640 -4581 -5616
rect -5949 -6960 -5925 -5640
rect -4605 -6960 -4581 -5640
rect -5949 -6984 -4581 -6960
rect -6743 -7081 -6423 -7039
rect -4245 -7039 -4203 -5561
rect -3967 -7039 -3925 -5561
rect -1747 -5561 -1427 -5519
rect -3451 -5640 -2083 -5616
rect -3451 -6960 -3427 -5640
rect -2107 -6960 -2083 -5640
rect -3451 -6984 -2083 -6960
rect -4245 -7081 -3925 -7039
rect -1747 -7039 -1705 -5561
rect -1469 -7039 -1427 -5561
rect 751 -5561 1071 -5519
rect -953 -5640 415 -5616
rect -953 -6960 -929 -5640
rect 391 -6960 415 -5640
rect -953 -6984 415 -6960
rect -1747 -7081 -1427 -7039
rect 751 -7039 793 -5561
rect 1029 -7039 1071 -5561
rect 3249 -5561 3569 -5519
rect 1545 -5640 2913 -5616
rect 1545 -6960 1569 -5640
rect 2889 -6960 2913 -5640
rect 1545 -6984 2913 -6960
rect 751 -7081 1071 -7039
rect 3249 -7039 3291 -5561
rect 3527 -7039 3569 -5561
rect 5747 -5561 6067 -5519
rect 4043 -5640 5411 -5616
rect 4043 -6960 4067 -5640
rect 5387 -6960 5411 -5640
rect 4043 -6984 5411 -6960
rect 3249 -7081 3569 -7039
rect 5747 -7039 5789 -5561
rect 6025 -7039 6067 -5561
rect 8245 -5561 8565 -5519
rect 6541 -5640 7909 -5616
rect 6541 -6960 6565 -5640
rect 7885 -6960 7909 -5640
rect 6541 -6984 7909 -6960
rect 5747 -7081 6067 -7039
rect 8245 -7039 8287 -5561
rect 8523 -7039 8565 -5561
rect 10743 -5561 11063 -5519
rect 9039 -5640 10407 -5616
rect 9039 -6960 9063 -5640
rect 10383 -6960 10407 -5640
rect 9039 -6984 10407 -6960
rect 8245 -7081 8565 -7039
rect 10743 -7039 10785 -5561
rect 11021 -7039 11063 -5561
rect 10743 -7081 11063 -7039
rect -9241 -7361 -8921 -7319
rect -10945 -7440 -9577 -7416
rect -10945 -8760 -10921 -7440
rect -9601 -8760 -9577 -7440
rect -10945 -8784 -9577 -8760
rect -9241 -8839 -9199 -7361
rect -8963 -8839 -8921 -7361
rect -6743 -7361 -6423 -7319
rect -8447 -7440 -7079 -7416
rect -8447 -8760 -8423 -7440
rect -7103 -8760 -7079 -7440
rect -8447 -8784 -7079 -8760
rect -9241 -8881 -8921 -8839
rect -6743 -8839 -6701 -7361
rect -6465 -8839 -6423 -7361
rect -4245 -7361 -3925 -7319
rect -5949 -7440 -4581 -7416
rect -5949 -8760 -5925 -7440
rect -4605 -8760 -4581 -7440
rect -5949 -8784 -4581 -8760
rect -6743 -8881 -6423 -8839
rect -4245 -8839 -4203 -7361
rect -3967 -8839 -3925 -7361
rect -1747 -7361 -1427 -7319
rect -3451 -7440 -2083 -7416
rect -3451 -8760 -3427 -7440
rect -2107 -8760 -2083 -7440
rect -3451 -8784 -2083 -8760
rect -4245 -8881 -3925 -8839
rect -1747 -8839 -1705 -7361
rect -1469 -8839 -1427 -7361
rect 751 -7361 1071 -7319
rect -953 -7440 415 -7416
rect -953 -8760 -929 -7440
rect 391 -8760 415 -7440
rect -953 -8784 415 -8760
rect -1747 -8881 -1427 -8839
rect 751 -8839 793 -7361
rect 1029 -8839 1071 -7361
rect 3249 -7361 3569 -7319
rect 1545 -7440 2913 -7416
rect 1545 -8760 1569 -7440
rect 2889 -8760 2913 -7440
rect 1545 -8784 2913 -8760
rect 751 -8881 1071 -8839
rect 3249 -8839 3291 -7361
rect 3527 -8839 3569 -7361
rect 5747 -7361 6067 -7319
rect 4043 -7440 5411 -7416
rect 4043 -8760 4067 -7440
rect 5387 -8760 5411 -7440
rect 4043 -8784 5411 -8760
rect 3249 -8881 3569 -8839
rect 5747 -8839 5789 -7361
rect 6025 -8839 6067 -7361
rect 8245 -7361 8565 -7319
rect 6541 -7440 7909 -7416
rect 6541 -8760 6565 -7440
rect 7885 -8760 7909 -7440
rect 6541 -8784 7909 -8760
rect 5747 -8881 6067 -8839
rect 8245 -8839 8287 -7361
rect 8523 -8839 8565 -7361
rect 10743 -7361 11063 -7319
rect 9039 -7440 10407 -7416
rect 9039 -8760 9063 -7440
rect 10383 -8760 10407 -7440
rect 9039 -8784 10407 -8760
rect 8245 -8881 8565 -8839
rect 10743 -8839 10785 -7361
rect 11021 -8839 11063 -7361
rect 10743 -8881 11063 -8839
<< properties >>
string FIXED_BBOX 8943 7320 10503 8880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 7.0 l 7.0 val 103.32 carea 2.00 cperi 0.19 nx 9 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
