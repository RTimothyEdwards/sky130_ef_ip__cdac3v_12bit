magic
tech sky130A
magscale 1 2
timestamp 1718247631
<< dnwell >>
rect 44121 -15586 48322 -14252
<< nwell >>
rect 44011 -14464 48431 -14149
rect 44011 -15380 46465 -14464
rect 48116 -15380 48431 -14464
rect 44011 -15695 48431 -15380
<< pwell >>
rect 46546 -15380 48116 -14464
<< psubdiff >>
rect 44052 -15873 44076 -15789
rect 48369 -15873 48393 -15789
<< mvpsubdiff >>
rect 46582 -14512 48080 -14500
rect 46582 -14546 46690 -14512
rect 46958 -14546 47116 -14512
rect 47542 -14546 47700 -14512
rect 47968 -14546 48080 -14512
rect 46582 -14558 48080 -14546
rect 46582 -14608 46640 -14558
rect 46582 -15236 46594 -14608
rect 46628 -15236 46640 -14608
rect 46582 -15286 46640 -15236
rect 47008 -14608 47066 -14558
rect 47008 -15236 47020 -14608
rect 47054 -15236 47066 -14608
rect 47008 -15286 47066 -15236
rect 47592 -14608 47650 -14558
rect 47592 -15236 47604 -14608
rect 47638 -15236 47650 -14608
rect 47592 -15286 47650 -15236
rect 48022 -14608 48080 -14558
rect 48022 -15236 48034 -14608
rect 48068 -15236 48080 -14608
rect 48022 -15286 48080 -15236
rect 46582 -15298 48080 -15286
rect 46582 -15332 46690 -15298
rect 46958 -15332 47116 -15298
rect 47542 -15332 47700 -15298
rect 47968 -15332 48080 -15298
rect 46582 -15344 48080 -15332
<< mvnsubdiff >>
rect 44078 -14235 48365 -14215
rect 44078 -14269 44158 -14235
rect 48285 -14269 48365 -14235
rect 44078 -14289 48365 -14269
rect 44078 -14295 44152 -14289
rect 44078 -15549 44098 -14295
rect 44132 -15549 44152 -14295
rect 48291 -14295 48365 -14289
rect 44273 -14514 46399 -14502
rect 44273 -14548 44381 -14514
rect 44807 -14548 44965 -14514
rect 45707 -14548 45865 -14514
rect 46291 -14548 46399 -14514
rect 44273 -14560 46399 -14548
rect 44273 -14610 44331 -14560
rect 44273 -15256 44285 -14610
rect 44319 -15256 44331 -14610
rect 44273 -15306 44331 -15256
rect 44857 -14610 44915 -14560
rect 44857 -15256 44869 -14610
rect 44903 -15256 44915 -14610
rect 44857 -15306 44915 -15256
rect 45757 -14610 45815 -14560
rect 45757 -15256 45769 -14610
rect 45803 -15256 45815 -14610
rect 45757 -15306 45815 -15256
rect 46341 -14610 46399 -14560
rect 46341 -15256 46353 -14610
rect 46387 -15256 46399 -14610
rect 46341 -15306 46399 -15256
rect 44273 -15318 46399 -15306
rect 44273 -15352 44381 -15318
rect 44807 -15352 44965 -15318
rect 45707 -15352 45865 -15318
rect 46291 -15352 46399 -15318
rect 44273 -15364 46399 -15352
rect 44078 -15555 44152 -15549
rect 48291 -15549 48311 -14295
rect 48345 -15549 48365 -14295
rect 48291 -15555 48365 -15549
rect 44078 -15575 48365 -15555
rect 44078 -15609 44158 -15575
rect 48285 -15609 48365 -15575
rect 44078 -15629 48365 -15609
<< psubdiffcont >>
rect 44076 -15873 48369 -15789
<< mvpsubdiffcont >>
rect 46690 -14546 46958 -14512
rect 47116 -14546 47542 -14512
rect 47700 -14546 47968 -14512
rect 46594 -15236 46628 -14608
rect 47020 -15236 47054 -14608
rect 47604 -15236 47638 -14608
rect 48034 -15236 48068 -14608
rect 46690 -15332 46958 -15298
rect 47116 -15332 47542 -15298
rect 47700 -15332 47968 -15298
<< mvnsubdiffcont >>
rect 44158 -14269 48285 -14235
rect 44098 -15549 44132 -14295
rect 44381 -14548 44807 -14514
rect 44965 -14548 45707 -14514
rect 45865 -14548 46291 -14514
rect 44285 -15256 44319 -14610
rect 44869 -15256 44903 -14610
rect 45769 -15256 45803 -14610
rect 46353 -15256 46387 -14610
rect 44381 -15352 44807 -15318
rect 44965 -15352 45707 -15318
rect 45865 -15352 46291 -15318
rect 48311 -15549 48345 -14295
rect 44158 -15609 48285 -15575
<< locali >>
rect 44098 -14269 44158 -14235
rect 48285 -14269 48345 -14235
rect 44098 -14295 48345 -14269
rect 44132 -14369 48311 -14295
rect 44132 -14514 44319 -14369
rect 46594 -14467 48101 -14449
rect 46594 -14504 46637 -14467
rect 47874 -14504 48101 -14467
rect 46594 -14512 48101 -14504
rect 44132 -14548 44381 -14514
rect 44807 -14548 44965 -14514
rect 45707 -14548 45865 -14514
rect 46291 -14548 46387 -14514
rect 44132 -14610 44319 -14548
rect 44132 -15256 44285 -14610
rect 44132 -15294 44319 -15256
rect 44869 -14610 44903 -14548
rect 44869 -15294 44903 -15256
rect 45769 -14610 45803 -14548
rect 45769 -15294 45803 -15256
rect 46353 -14610 46387 -14548
rect 46353 -15294 46387 -15256
rect 46594 -14546 46690 -14512
rect 46958 -14546 47116 -14512
rect 47542 -14546 47700 -14512
rect 47968 -14546 48101 -14512
rect 46594 -14566 48101 -14546
rect 46594 -14608 46628 -14566
rect 44132 -15318 46388 -15294
rect 44132 -15352 44381 -15318
rect 44807 -15345 44965 -15318
rect 45707 -15345 45865 -15318
rect 46291 -15345 46388 -15318
rect 44132 -15380 44500 -15352
rect 46363 -15380 46388 -15345
rect 44132 -15388 46388 -15380
rect 46594 -15298 46628 -15236
rect 47020 -14608 47054 -14566
rect 47020 -15298 47054 -15236
rect 47604 -14608 47638 -14566
rect 47604 -15298 47638 -15236
rect 48034 -14608 48068 -14566
rect 48034 -15298 48068 -15236
rect 46594 -15332 46690 -15298
rect 46958 -15332 47116 -15298
rect 47542 -15332 47700 -15298
rect 47968 -15332 48068 -15298
rect 46594 -15355 48066 -15332
rect 44132 -15473 44319 -15388
rect 46594 -15401 46616 -15355
rect 48048 -15401 48066 -15355
rect 46594 -15411 48066 -15401
rect 48160 -15473 48311 -14369
rect 44132 -15549 48311 -15473
rect 44098 -15575 48345 -15549
rect 44098 -15609 44158 -15575
rect 48285 -15609 48345 -15575
rect 46757 -15736 47157 -15714
rect 46757 -15789 46778 -15736
rect 47140 -15789 47157 -15736
rect 44060 -15873 44076 -15789
rect 48369 -15873 48385 -15789
rect 46757 -15935 46778 -15873
rect 47140 -15935 47157 -15873
rect 46757 -15952 47157 -15935
<< viali >>
rect 46637 -14504 47874 -14467
rect 44500 -15352 44807 -15345
rect 44807 -15352 44965 -15345
rect 44965 -15352 45707 -15345
rect 45707 -15352 45865 -15345
rect 45865 -15352 46291 -15345
rect 46291 -15352 46363 -15345
rect 44500 -15380 46363 -15352
rect 46616 -15401 48048 -15355
rect 46778 -15789 47140 -15736
rect 45020 -15873 45210 -15789
rect 46778 -15873 47140 -15789
rect 46778 -15935 47140 -15873
<< metal1 >>
rect 44011 -14426 48101 -14409
rect 44011 -14543 45575 -14426
rect 45942 -14467 48101 -14426
rect 45942 -14504 46637 -14467
rect 47874 -14504 48101 -14467
rect 45942 -14543 48101 -14504
rect 44011 -14555 48101 -14543
rect 44011 -15325 46402 -15311
rect 44011 -15345 44973 -15325
rect 45341 -15345 46402 -15325
rect 44011 -15380 44500 -15345
rect 46363 -15380 46402 -15345
rect 44011 -15444 44973 -15380
rect 45341 -15444 46402 -15380
rect 44011 -15457 46402 -15444
rect 46594 -15355 48119 -15311
rect 46594 -15401 46616 -15355
rect 48048 -15401 48119 -15355
rect 46594 -15457 48119 -15401
rect 46757 -15736 47157 -15714
rect 45007 -15789 45224 -15779
rect 45007 -15873 45020 -15789
rect 45210 -15873 45224 -15789
rect 45007 -15884 45224 -15873
rect 46757 -15935 46778 -15736
rect 47140 -15935 47157 -15736
rect 46757 -15952 47157 -15935
<< via1 >>
rect 45575 -14543 45942 -14426
rect 44973 -15345 45341 -15325
rect 44973 -15380 45341 -15345
rect 44973 -15444 45341 -15380
rect 46778 -15935 47140 -15736
<< metal2 >>
rect 45557 -14336 45957 -14318
rect 45557 -14543 45574 -14336
rect 45942 -14543 45957 -14336
rect 45557 -14555 45957 -14543
rect 44957 -15325 45357 -15311
rect 44957 -15512 44973 -15325
rect 45342 -15512 45357 -15325
rect 44957 -15525 45357 -15512
rect 46757 -15736 47157 -15714
rect 46757 -15935 46778 -15736
rect 47140 -15935 47157 -15736
rect 46757 -15952 47157 -15935
<< via2 >>
rect 45574 -14426 45942 -14336
rect 45574 -14543 45575 -14426
rect 45575 -14543 45942 -14426
rect 44973 -15444 45341 -15325
rect 45341 -15444 45342 -15325
rect 44973 -15512 45342 -15444
rect 46778 -15935 47140 -15736
<< metal3 >>
rect 45557 -14336 45957 -14318
rect 45557 -14543 45574 -14336
rect 45942 -14543 45957 -14336
rect 45557 -14555 45957 -14543
rect 44957 -15325 45357 -15311
rect 44957 -15512 44973 -15325
rect 45342 -15512 45357 -15325
rect 44957 -15525 45357 -15512
rect 46757 -15736 47157 -15714
rect 46757 -15935 46778 -15736
rect 47140 -15935 47157 -15736
rect 46757 -15952 47157 -15935
<< labels >>
flabel metal1 44011 -14555 44167 -14409 0 FreeSans 800 0 0 0 avss
port 5 nsew
flabel metal1 44011 -15457 44167 -15311 0 FreeSans 800 0 0 0 avdd
port 4 nsew
<< end >>
