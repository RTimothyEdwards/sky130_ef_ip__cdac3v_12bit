magic
tech sky130A
magscale 1 2
timestamp 1722784074
<< metal3 >>
rect 81341 -31719 81401 -31579
rect 81031 -32029 82511 -31719
rect 81031 -32089 82651 -32029
rect 81031 -32840 82511 -32089
rect 80891 -32900 82511 -32840
rect 81031 -33210 82511 -32900
rect 82141 -33350 82201 -33210
<< mimcap >>
rect 81071 -31799 82471 -31759
rect 81071 -33130 81111 -31799
rect 82431 -33130 82471 -31799
rect 81071 -33170 82471 -33130
<< mimcapcontact >>
rect 81111 -33130 82431 -31799
<< metal4 >>
rect 81741 -31679 81801 -31579
rect 80991 -31799 82551 -31679
rect 80991 -32434 81111 -31799
rect 80891 -32494 81111 -32434
rect 80991 -33130 81111 -32494
rect 82431 -32434 82551 -31799
rect 82431 -32494 82651 -32434
rect 82431 -33130 82551 -32494
rect 80991 -33250 82551 -33130
rect 81741 -33350 81801 -33250
<< mimcap2 >>
rect 81071 -31799 82471 -31759
rect 81071 -33130 81111 -31799
rect 82431 -33130 82471 -31799
rect 81071 -33170 82471 -33130
<< mimcap2contact >>
rect 81111 -33130 82431 -31799
<< metal5 >>
rect 82011 -31775 82331 -31084
rect 81087 -31799 82455 -31775
rect 81087 -31899 81111 -31799
rect 80396 -32219 81111 -31899
rect 81087 -33130 81111 -32219
rect 82431 -32710 82455 -31799
rect 82431 -33030 83146 -32710
rect 82431 -33130 82455 -33030
rect 81087 -33154 82455 -33130
rect 81211 -33846 81531 -33154
<< properties >>
string cdac_ratioed_cap gencell
<< end >>
