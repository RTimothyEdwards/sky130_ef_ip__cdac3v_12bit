magic
tech sky130A
magscale 1 2
timestamp 1718247631
<< error_s >>
rect 1876 4154 2249 4159
rect 1876 3945 1881 4154
rect 2244 3945 2249 4154
rect 1876 3940 2249 3945
rect 1877 3514 2245 3519
rect 1877 3360 1882 3514
rect 2240 3360 2245 3514
rect 1877 3355 2245 3360
rect 1275 3159 1654 3164
rect 1275 2961 1277 3159
rect 1649 2961 1654 3159
rect 1275 2956 1654 2961
rect 3083 2742 3445 2747
rect 3083 2561 3088 2742
rect 3440 2561 3445 2742
rect 3083 2556 3445 2561
rect 2476 1840 2848 1845
rect 2476 1701 2481 1840
rect 2843 1701 2848 1840
rect 2476 1696 2848 1701
rect 3075 839 3453 844
rect 3075 619 3080 839
rect 3448 619 3453 839
rect 3075 614 3453 619
rect 2477 -254 2853 -249
rect 2477 -358 2482 -254
rect 2848 -358 2853 -254
rect 2477 -363 2853 -358
rect 3082 -1104 3446 -1099
rect 3082 -1287 3087 -1104
rect 3441 -1287 3446 -1104
rect 3082 -1292 3446 -1287
rect 1275 -1507 1649 -1502
rect 1275 -1697 1280 -1507
rect 1644 -1697 1649 -1507
rect 1275 -1702 1649 -1697
rect 1876 -1904 2244 -1899
rect 1876 -2058 1881 -1904
rect 2239 -2058 2244 -1904
rect 1876 -2063 2244 -2058
rect 1874 -2488 2249 -2483
rect 1874 -2675 1879 -2488
rect 2244 -2675 2249 -2488
rect 1874 -2680 2249 -2675
<< viali >>
rect 3083 2556 3445 2747
rect 3082 -1292 3446 -1099
<< metal1 >>
rect 1272 3104 1276 3164
rect 3064 2747 3464 2765
rect 3064 2556 3083 2747
rect 3445 2556 3464 2747
rect 3064 2538 3464 2556
rect 721 2096 783 2103
rect 721 1976 726 2096
rect 778 1976 783 2096
rect 721 1969 783 1976
rect 418 1418 809 1668
rect 318 630 518 830
rect 319 -438 519 -238
rect 721 -516 783 -509
rect 721 -635 726 -516
rect 778 -635 783 -516
rect 721 -643 783 -635
rect 320 -946 520 -746
rect 3064 -1099 3464 -1082
rect 3064 -1292 3082 -1099
rect 3446 -1292 3464 -1099
rect 3064 -1312 3464 -1292
rect 817 -2616 1017 -2470
<< via1 >>
rect 1876 3939 2249 4058
rect 1276 3104 1656 3164
rect 3083 2556 3445 2747
rect 726 1976 778 2096
rect 2476 1696 2848 1753
rect 3075 614 3453 844
rect 2477 -295 2854 -238
rect 726 -635 778 -516
rect 3082 -1292 3446 -1099
rect 1274 -1706 1650 -1637
rect 1874 -2602 2249 -2483
<< metal2 >>
rect 1863 4159 2264 4180
rect 1863 3939 1876 4159
rect 2249 3939 2264 4159
rect 1863 3928 2264 3939
rect 4734 3573 4934 3773
rect 1264 3164 1664 3172
rect 1264 2956 1275 3164
rect 1656 3104 1664 3164
rect 1654 2956 1664 3104
rect 1264 2945 1664 2956
rect 3064 2747 3464 2765
rect 3064 2556 3083 2747
rect 3445 2556 3464 2747
rect 3064 2538 3464 2556
rect 721 2096 783 2103
rect 721 1976 726 2096
rect 778 1976 783 2096
rect 721 1969 783 1976
rect 721 -509 759 1969
rect 2464 1845 2864 1857
rect 2464 1696 2476 1845
rect 2848 1696 2864 1845
rect 3064 844 3464 854
rect 3064 614 3075 844
rect 3453 614 3464 844
rect 3064 604 3464 614
rect 2464 -238 2864 -237
rect 2464 -363 2477 -238
rect 2854 -295 2864 -238
rect 2853 -363 2864 -295
rect 2464 -376 2864 -363
rect 721 -516 783 -509
rect 721 -635 726 -516
rect 778 -635 783 -516
rect 721 -643 783 -635
rect 3064 -1099 3464 -1082
rect 3064 -1292 3082 -1099
rect 3446 -1292 3464 -1099
rect 3064 -1312 3464 -1292
rect 1264 -1502 1664 -1489
rect 1264 -1637 1275 -1502
rect 1649 -1637 1664 -1502
rect 1264 -1706 1274 -1637
rect 1650 -1706 1664 -1637
rect 1264 -1714 1664 -1706
rect 4734 -2316 4934 -2116
rect 1864 -2483 2264 -2470
rect 1864 -2680 1874 -2483
rect 2249 -2680 2264 -2483
rect 1864 -2698 2264 -2680
<< via2 >>
rect 1876 4058 2249 4159
rect 1876 3940 2249 4058
rect 1877 3355 2245 3519
rect 1275 3104 1276 3164
rect 1276 3104 1654 3164
rect 1275 2956 1654 3104
rect 3083 2556 3445 2747
rect 2476 1753 2848 1845
rect 2476 1696 2848 1753
rect 3075 614 3453 844
rect 2477 -295 2853 -249
rect 2477 -363 2853 -295
rect 3082 -1292 3446 -1099
rect 1275 -1637 1649 -1502
rect 1275 -1702 1649 -1637
rect 1876 -2063 2244 -1899
rect 1874 -2602 2249 -2483
rect 1874 -2680 2249 -2602
<< metal3 >>
rect 1272 2956 1275 3164
use simple_analog_switch_ena1v8  simple_analog_switch_ena1v8_0 ../../../dependencies/sky130_ef_ip__analog_switches/mag
timestamp 1718247631
transform 1 0 318 0 -1 4334
box 0 0 4420 3648
use simple_analog_switch_ena1v8  simple_analog_switch_ena1v8_1
timestamp 1718247631
transform 1 0 318 0 1 -2876
box 0 0 4420 3648
<< labels >>
flabel metal1 320 -946 520 -746 0 FreeSans 256 0 0 0 RST
port 5 nsew
flabel metal1 318 630 518 830 0 FreeSans 256 0 0 0 DVSS
port 6 nsew
flabel metal1 319 -438 519 -238 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal1 443 1442 643 1642 0 FreeSans 256 0 0 0 AVDD
port 2 nsew
flabel metal1 817 -2616 1017 -2470 0 FreeSans 256 0 0 0 AVSS
port 4 nsew
flabel metal2 4734 3573 4934 3773 0 FreeSans 256 0 0 0 VP2
port 1 nsew
flabel metal2 4734 -2316 4934 -2116 0 FreeSans 256 0 0 0 VP1
port 0 nsew
<< end >>
