magic
tech sky130A
magscale 1 2
timestamp 1731116683
<< dnwell >>
rect 53466 -9213 56720 -8556
rect 85693 -9164 88946 -8556
rect 53510 -9306 56764 -9213
rect 84771 -10934 88972 -10498
rect 53467 -12960 56720 -12238
rect 85693 -12960 88946 -12268
<< nwell >>
rect 85584 -9061 89055 -8560
rect 84662 -10825 89082 -10607
rect 53359 -13008 56830 -12813
rect 85583 -12953 89054 -12371
<< viali >>
rect 58720 12899 83690 12933
rect 58631 -34472 58665 12845
rect 83747 -34470 83781 12837
rect 58722 -34559 83692 -34525
<< metal1 >>
rect 87993 14759 88037 14793
rect 87993 14660 88037 14691
rect 57694 13813 57706 13826
rect 57681 13765 57706 13813
rect 57925 13813 57937 13826
rect 84498 13816 84508 13820
rect 81689 13813 84508 13816
rect 57925 13768 84508 13813
rect 84674 13768 84683 13820
rect 57925 13765 82020 13768
rect 53335 13669 71029 13717
rect 73635 13669 89082 13717
rect 53239 13573 61188 13621
rect 63475 13573 89177 13621
rect 53142 13477 66185 13525
rect 68465 13477 89273 13525
rect 53046 13381 80253 13429
rect 80925 13381 89368 13429
rect 80205 13333 80253 13381
rect 52949 13285 75727 13333
rect 75994 13285 80108 13333
rect 80205 13285 83639 13333
rect 84364 13285 89464 13333
rect 75679 13237 75727 13285
rect 80059 13239 80107 13285
rect 84364 13239 84456 13285
rect 52849 13189 75605 13237
rect 75679 13189 78562 13237
rect 80059 13191 84456 13239
rect 88767 13189 89562 13237
rect 75557 13145 75605 13189
rect 52856 10694 53466 10742
rect 52952 3490 53506 3538
rect 53048 -3715 53453 -3667
rect 56963 -8434 57004 13133
rect 53593 -8475 57004 -8434
rect 57048 -8528 57089 13133
rect 75557 13097 88636 13145
rect 88767 13045 88815 13189
rect 85980 12997 88815 13045
rect 58611 12933 83801 12953
rect 58611 12899 58720 12933
rect 83690 12899 83801 12933
rect 58611 12879 83801 12899
rect 58611 12845 58685 12879
rect 53503 -8569 57089 -8528
rect 53089 -15323 53462 -15275
rect 53089 -22526 53456 -22478
rect 53089 -29732 53501 -29672
rect 58611 -34472 58631 12845
rect 58665 -34472 58685 12845
rect 58611 -34505 58685 -34472
rect 83727 12837 83801 12879
rect 83727 -34470 83747 12837
rect 83781 -34470 83801 12837
rect 88909 10698 89507 10741
rect 88909 10693 89557 10698
rect 88933 3490 89469 3538
rect 88931 -3714 89372 -3666
rect 88922 -15322 89306 -15274
rect 88958 -22526 89322 -22478
rect 88912 -29734 89329 -29661
rect 83727 -34505 83801 -34470
rect 58611 -34525 83801 -34505
rect 58611 -34559 58722 -34525
rect 83692 -34559 83801 -34525
rect 58611 -34579 83801 -34559
rect 58611 -34690 58685 -34579
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -34948 58685 -34939
rect 83727 -34698 83801 -34579
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 83727 -34955 83801 -34947
<< via1 >>
rect 67193 15465 68325 15613
rect 74728 14929 75860 15002
rect 53998 14659 54340 14894
rect 88037 14660 88414 14890
rect 67192 13939 68325 14087
rect 57706 13765 57925 13826
rect 84508 13768 84674 13820
rect 57778 12794 57854 12980
rect 84559 12794 84635 12977
rect 58619 -34939 58678 -34690
rect 83734 -34947 83793 -34698
<< metal2 >>
rect 54231 15270 54431 15691
rect 56731 15278 56931 15691
rect 59240 15258 59440 15689
rect 61738 15269 61938 15686
rect 64226 15272 64426 15683
rect 66724 15269 66924 15678
rect 67192 15613 68325 15674
rect 67192 15465 67193 15613
rect 53989 14894 54350 14901
rect 53989 14659 53998 14894
rect 54340 14659 54350 14894
rect 53989 14651 54350 14659
rect 67192 14087 68325 15465
rect 69204 15277 69404 15673
rect 71707 15264 71907 15681
rect 74204 15267 74404 15673
rect 52859 10690 52907 13362
rect 52955 3485 53003 13445
rect 53051 -3719 53099 13549
rect 53147 -15369 53195 13650
rect 53243 -22539 53291 13747
rect 53339 -29684 53387 13824
rect 53627 13805 53663 13983
rect 56057 13878 56093 13947
rect 56057 13842 57083 13878
rect 58537 13859 58605 13989
rect 53627 13769 57000 13805
rect 56964 13114 57000 13769
rect 57047 13118 57083 13842
rect 57783 13826 58605 13859
rect 57694 13765 57706 13826
rect 57925 13791 58605 13826
rect 57925 13765 57937 13791
rect 57783 12986 57851 13765
rect 61047 13580 61091 13960
rect 63543 13596 63587 13960
rect 66039 13492 66083 13960
rect 74728 15002 75860 15672
rect 76712 15261 76912 15677
rect 79201 15260 79401 15680
rect 81703 15255 81903 15678
rect 84207 15264 84407 15683
rect 86689 15259 86889 15678
rect 74728 14497 75860 14929
rect 88024 14890 88424 14901
rect 88024 14660 88037 14890
rect 88414 14660 88424 14890
rect 88024 14651 88424 14660
rect 74728 14149 74753 14497
rect 75837 14149 75860 14497
rect 67192 13924 68325 13939
rect 67192 13577 67221 13924
rect 68291 13577 68325 13924
rect 67192 13552 68325 13577
rect 68535 13496 68579 13960
rect 71031 13691 71075 13964
rect 73527 13839 73571 13960
rect 73527 13795 73573 13839
rect 73529 13691 73573 13795
rect 74728 13714 75860 14149
rect 76023 13295 76067 13960
rect 78519 13195 78563 13960
rect 81015 13413 81059 13960
rect 83511 13308 83555 13960
rect 84498 13768 84508 13820
rect 84674 13768 84685 13820
rect 84565 12986 84629 13768
rect 86007 13003 86051 13960
rect 88503 13116 88547 13963
rect 57778 12980 57854 12986
rect 57778 12786 57854 12794
rect 84559 12977 84635 12986
rect 84559 12786 84635 12794
rect 53462 -10689 53500 -8524
rect 53551 -10485 53589 -8428
rect 57595 -9382 57659 -9322
rect 57595 -9823 57659 -9664
rect 53551 -10523 53730 -10485
rect 53692 -10705 53730 -10523
rect 53543 -10743 53730 -10705
rect 53543 -10840 53581 -10743
rect 57595 -11967 57659 -11601
rect 57595 -12288 57659 -12249
rect 89029 -29735 89077 13849
rect 89125 -22535 89173 13742
rect 89221 -15347 89269 13661
rect 89317 -3749 89365 13564
rect 89413 3485 89461 13478
rect 89509 10895 89557 13371
rect 89509 10686 89557 10698
rect 58611 -34690 58685 -34682
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -36047 58685 -34939
rect 83727 -34698 83801 -34690
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 68751 -35460 70341 -35417
rect 68751 -35798 68783 -35460
rect 70303 -35798 70341 -35460
rect 58611 -36058 58735 -36047
rect 58611 -36434 58624 -36058
rect 58724 -36434 58735 -36058
rect 58611 -36441 58735 -36434
rect 58612 -36446 58735 -36441
rect 68751 -36556 70341 -35798
rect 72201 -36081 73791 -36042
rect 83727 -36047 83801 -34947
rect 72201 -36419 72237 -36081
rect 73757 -36419 73791 -36081
rect 72201 -36568 73791 -36419
rect 83672 -36059 83801 -36047
rect 83672 -36435 83686 -36059
rect 83789 -36435 83801 -36059
rect 83672 -36447 83801 -36435
<< via2 >>
rect 53998 14659 54340 14894
rect 88037 14660 88414 14890
rect 74753 14149 75837 14497
rect 67221 13577 68291 13924
rect 57595 -9664 57659 -9382
rect 57595 -12249 57659 -11967
rect 68783 -35798 70303 -35460
rect 58624 -36434 58724 -36058
rect 72237 -36419 73757 -36081
rect 83686 -36435 83789 -36059
<< metal3 >>
rect 53989 14894 54389 14942
rect 53989 14659 53998 14894
rect 54340 14659 54389 14894
rect 53989 13063 54389 14659
rect 88024 14890 88424 14927
rect 88024 14660 88037 14890
rect 88414 14660 88424 14890
rect 74753 14497 75837 14498
rect 65040 14202 65240 14402
rect 64616 13678 64816 13878
rect 88024 13066 88424 14660
rect 57444 10300 57452 10364
rect 57681 10300 58425 10364
rect 84059 10176 85266 10240
rect 57134 7820 58405 7884
rect 57146 2736 58413 2800
rect 83551 2736 84399 2800
rect 84606 2736 84613 2800
rect 83933 256 85271 320
rect 57134 -4704 58320 -4640
rect 83918 -7060 85398 -6996
rect 57590 -9382 57664 -9376
rect 57590 -9664 57595 -9382
rect 57659 -9600 57664 -9382
rect 89066 -9592 89295 -9586
rect 84666 -9600 84873 -9594
rect 57659 -9664 58900 -9600
rect 83980 -9664 84671 -9600
rect 84867 -9664 84873 -9600
rect 57590 -9669 57664 -9664
rect 84666 -9670 84873 -9664
rect 89066 -9667 89075 -9592
rect 89286 -9600 89295 -9592
rect 89380 -9600 89580 -9514
rect 89286 -9664 89580 -9600
rect 89286 -9667 89295 -9664
rect 89066 -9674 89295 -9667
rect 89380 -9714 89580 -9664
rect 53096 -10372 53248 -10362
rect 53096 -10781 53108 -10372
rect 53237 -10781 53248 -10372
rect 53096 -10794 53248 -10781
rect 53096 -11173 53247 -10794
rect 57590 -11967 57664 -11962
rect 57590 -12249 57595 -11967
rect 57659 -12031 58919 -11967
rect 57659 -12249 57664 -12031
rect 83840 -12036 84037 -11972
rect 57590 -12255 57664 -12249
rect 57014 -14635 58370 -14571
rect 83950 -16991 85256 -16927
rect 57162 -21951 58447 -21887
rect 53226 -24291 53363 -24278
rect 53226 -24333 53243 -24291
rect 53077 -24468 53243 -24333
rect 53226 -24685 53243 -24468
rect 53349 -24685 53363 -24291
rect 54633 -24475 55033 -24319
rect 58042 -24363 58280 -24351
rect 58042 -24429 58054 -24363
rect 58266 -24367 58280 -24363
rect 58266 -24429 58410 -24367
rect 58042 -24431 58410 -24429
rect 83988 -24431 85276 -24367
rect 58042 -24445 58280 -24431
rect 53226 -24704 53363 -24685
rect 83963 -29515 85267 -29451
rect 54633 -31901 55033 -31860
rect 57141 -31871 58330 -31807
rect 54633 -32023 54649 -31901
rect 55017 -32023 55033 -31901
rect 54633 -32057 55033 -32023
rect 58042 -31943 58816 -31931
rect 58042 -32009 58054 -31943
rect 58266 -31995 58816 -31943
rect 83980 -31995 84409 -31931
rect 84644 -31995 84651 -31931
rect 58266 -32009 58280 -31995
rect 58042 -32025 58280 -32009
rect 70215 -34911 70415 -34711
rect 53497 -35185 53696 -34986
rect 70614 -35211 70814 -35011
rect 65838 -35733 66038 -35533
rect 65303 -36348 65503 -36148
<< via3 >>
rect 54595 10276 54983 10399
rect 57452 10300 57681 10364
rect 84399 2736 84606 2800
rect 87436 2703 87813 2834
rect 84671 -9664 84867 -9600
rect 89075 -9667 89286 -9592
rect 53108 -10781 53237 -10372
rect 56986 -10947 57151 -10416
rect 53243 -24685 53349 -24291
rect 58054 -24429 58266 -24363
rect 54649 -32023 55017 -31901
rect 58054 -32009 58266 -31943
rect 84409 -31995 84644 -31931
rect 87430 -32014 87818 -31910
<< metal4 >>
rect 54589 10399 54989 10400
rect 54589 10276 54595 10399
rect 54983 10364 54989 10399
rect 57451 10364 57682 10365
rect 54983 10300 57452 10364
rect 57681 10300 57682 10364
rect 54983 10276 54989 10300
rect 57451 10299 57682 10300
rect 54589 10275 54989 10276
rect 87424 2834 87824 2845
rect 84398 2800 84607 2801
rect 87424 2800 87436 2834
rect 84398 2736 84399 2800
rect 84606 2736 87436 2800
rect 84398 2735 84607 2736
rect 87424 2703 87436 2736
rect 87813 2703 87824 2834
rect 87424 2691 87824 2703
rect 89066 -9592 89295 -9586
rect 84666 -9600 84873 -9594
rect 89066 -9600 89075 -9592
rect 84666 -9664 84671 -9600
rect 84867 -9664 89075 -9600
rect 84666 -9670 84873 -9664
rect 89066 -9667 89075 -9664
rect 89286 -9667 89295 -9592
rect 89066 -9674 89295 -9667
rect 53096 -10372 53248 -10362
rect 53096 -10781 53108 -10372
rect 53237 -10622 53248 -10372
rect 56970 -10416 57166 -10401
rect 56970 -10622 56986 -10416
rect 53237 -10774 56986 -10622
rect 53237 -10781 53248 -10774
rect 53096 -10794 53248 -10781
rect 56970 -10947 56986 -10774
rect 57151 -10947 57166 -10416
rect 56970 -10965 57166 -10947
rect 53226 -24291 53363 -24278
rect 53226 -24685 53243 -24291
rect 53349 -24369 53363 -24291
rect 58042 -24363 58280 -24351
rect 58042 -24369 58054 -24363
rect 53349 -24429 58054 -24369
rect 58266 -24429 58280 -24363
rect 53349 -24685 53363 -24429
rect 58042 -24445 58280 -24429
rect 53226 -24704 53363 -24685
rect 54631 -31901 55037 -31883
rect 54631 -32023 54649 -31901
rect 55017 -31933 55037 -31901
rect 87424 -31910 87824 -31909
rect 84408 -31931 84645 -31930
rect 87424 -31931 87430 -31910
rect 58042 -31933 58280 -31931
rect 55017 -31943 58280 -31933
rect 55017 -31993 58054 -31943
rect 55017 -32023 55037 -31993
rect 54631 -32039 55037 -32023
rect 58042 -32009 58054 -31993
rect 58266 -32009 58280 -31943
rect 84408 -31995 84409 -31931
rect 84644 -31995 87430 -31931
rect 84408 -31996 84645 -31995
rect 58042 -32025 58280 -32009
rect 87424 -32014 87430 -31995
rect 87818 -32014 87824 -31910
rect 87424 -32015 87824 -32014
use cdac_dummy_switch  cdac_dummy_switch_1
timestamp 1731099133
transform -1 0 133093 0 1 5088
box 44011 -15952 48431 -14149
use cdac_dummy_switch  cdac_dummy_switch_2
timestamp 1731099133
transform -1 0 133093 0 -1 -26520
box 44011 -15952 48431 -14149
use cdac_lvlshift_array  cdac_lvlshift_array_0
timestamp 1731114850
transform 1 0 -395 0 1 -788
box 53822 14704 89378 16424
use cdac_via_3cut  cdac_via_3cut_0
timestamp 1718247631
transform 1 0 708 0 1 36628
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_1
timestamp 1718247631
transform 1 0 709 0 1 3409
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_2
timestamp 1718247631
transform 1 0 708 0 1 10604
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_3
timestamp 1718247631
transform 1 0 708 0 1 17763
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_4
timestamp 1718247631
transform 1 0 709 0 1 29419
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_5
timestamp 1718247631
transform 1 0 36175 0 1 17813
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_6
timestamp 1718247631
transform 1 0 705 0 1 43828
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_7
timestamp 1718247631
transform 1 0 36172 0 1 3404
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_8
timestamp 1718247631
transform 1 0 36176 0 1 10609
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_9
timestamp 1718247631
transform 1 0 36167 0 1 29422
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_10
timestamp 1718247631
transform 1 0 36182 0 1 43834
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_11
timestamp 1718247631
transform 1 0 36176 0 1 36626
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_12
timestamp 1718247631
transform -1 0 106247 0 -1 -41658
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_13
timestamp 1718247631
transform 1 0 213 0 1 46421
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_14
timestamp 1718247631
transform 1 0 308 0 1 46517
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_15
timestamp 1718247631
transform 1 0 404 0 1 46613
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_16
timestamp 1718247631
transform 1 0 501 0 1 46708
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_17
timestamp 1718247631
transform 1 0 595 0 1 46803
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_18
timestamp 1718247631
transform 1 0 36768 0 1 46325
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_19
timestamp 1718247631
transform 1 0 36670 0 1 46419
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_20
timestamp 1718247631
transform 1 0 36574 0 1 46517
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_21
timestamp 1718247631
transform 1 0 36478 0 1 46612
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_22
timestamp 1718247631
transform 1 0 36381 0 1 46709
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_23
timestamp 1718247631
transform 1 0 36286 0 1 46805
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_24
timestamp 1718247631
transform 0 1 104033 -1 0 66458
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_25
timestamp 1718247631
transform 0 1 94111 -1 0 66359
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_26
timestamp 1718247631
transform 0 1 106653 -1 0 66463
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_27
timestamp 1718247631
transform 0 1 99107 -1 0 66269
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_28
timestamp 1718247631
transform 0 1 96603 -1 0 66364
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_29
timestamp 1718247631
transform 0 1 101602 -1 0 66269
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_30
timestamp 1718247631
transform 0 1 111586 -1 0 65977
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_31
timestamp 1718247631
transform 0 1 116593 -1 0 66081
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_32
timestamp 1718247631
transform 0 1 114058 -1 0 66173
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_33
timestamp 1718247631
transform 0 1 109128 -1 0 66070
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_34
timestamp 1718247631
transform 0 1 119100 -1 0 65788
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_35
timestamp 1718247631
transform 0 1 121568 -1 0 65887
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_36
timestamp 1718247631
transform 1 0 116 0 1 43829
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_38
timestamp 1718247631
transform 1 0 212 0 1 36624
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_39
timestamp 1718247631
transform 1 0 308 0 1 29419
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_40
timestamp 1718247631
transform 1 0 405 0 1 17763
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_41
timestamp 1718247631
transform 1 0 501 0 1 10604
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_42
timestamp 1718247631
transform 1 0 597 0 1 3406
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_43
timestamp 1718247631
transform 1 0 36767 0 1 43829
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_44
timestamp 1718247631
transform 1 0 36670 0 1 36626
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_45
timestamp 1718247631
transform 1 0 36571 0 1 29422
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_46
timestamp 1718247631
transform 1 0 36481 0 1 17812
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_47
timestamp 1718247631
transform 1 0 36382 0 1 10606
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_48
timestamp 1718247631
transform 1 0 36286 0 1 3404
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_49
timestamp 1718247631
transform 1 0 4303 0 1 46075
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_50
timestamp 1718247631
transform 1 0 4219 0 1 46073
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_51
timestamp 1718247631
transform 1 0 116 0 1 46324
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_52
timestamp 1718247631
transform 0 1 86685 -1 0 44315
box 52740 -33138 52792 -32927
use EF_SW_RST  x1
timestamp 1731116066
transform 1 0 52725 0 -1 -9897
box 563 -2876 4983 4338
use EF_AMUX0201_ARRAY1  x3
timestamp 1731116499
transform 0 1 62083 -1 0 14841
box 320 -8725 51288 26972
use EF_BANK_CAP_12  x4
timestamp 1731114039
transform 1 0 0 0 1 -8000
box 58243 -26640 84124 21013
<< labels >>
flabel metal3 64616 13678 64816 13878 0 FreeSans 256 90 0 0 DVSS
port 12 nsew
flabel metal3 65040 14202 65240 14402 0 FreeSans 256 90 0 0 DVDD
port 11 nsew
flabel metal3 83840 -12036 84037 -11972 0 FreeSans 480 0 0 0 OUTNC
port 22 nsew
flabel metal3 53077 -24468 53216 -24333 0 FreeSans 480 0 0 0 Vref
port 25 nsew
flabel metal2 56731 15491 56931 15691 0 FreeSans 480 0 0 0 RST
port 17 nsew
flabel metal2 54231 15507 54431 15691 0 FreeSans 480 0 0 0 HOLD
port 27 nsew
flabel metal2 59240 15489 59440 15689 0 FreeSans 480 0 0 0 SELD0
port 23 nsew
flabel metal2 61738 15486 61938 15686 0 FreeSans 480 0 0 0 SELD1
port 24 nsew
flabel metal2 64226 15483 64426 15683 0 FreeSans 480 0 0 0 SELD2
port 2 nsew
flabel metal2 66724 15478 66924 15678 0 FreeSans 480 0 0 0 SELD3
port 3 nsew
flabel metal2 69204 15473 69404 15673 0 FreeSans 480 0 0 0 SELD4
port 4 nsew
flabel metal2 71707 15481 71907 15681 0 FreeSans 480 0 0 0 SELD5
port 5 nsew
flabel metal2 74204 15473 74404 15673 0 FreeSans 480 0 0 0 SELD6
port 6 nsew
flabel metal2 76712 15477 76912 15677 0 FreeSans 480 0 0 0 SELD7
port 7 nsew
flabel metal2 79201 15480 79401 15680 0 FreeSans 480 0 0 0 SELD8
port 8 nsew
flabel metal2 86689 15478 86889 15678 0 FreeSans 480 0 0 0 SELD11
port 21 nsew
flabel metal2 84207 15483 84407 15683 0 FreeSans 480 0 0 0 SELD10
port 19 nsew
flabel metal2 81703 15478 81903 15678 0 FreeSans 480 0 0 0 SELD9
port 9 nsew
flabel metal3 70614 -35211 70814 -35011 0 FreeSans 256 90 0 0 VH
port 14 nsew
flabel metal3 70215 -34911 70415 -34711 0 FreeSans 256 90 0 0 VL
port 15 nsew
flabel metal3 65303 -36348 65503 -36148 0 FreeSans 256 90 0 0 VDD
port 10 nsew
flabel metal3 65838 -35733 66038 -35533 0 FreeSans 256 90 0 0 VSS
port 13 nsew
flabel metal3 89380 -9714 89580 -9514 0 FreeSans 480 0 0 0 OUT
port 16 nsew
flabel metal3 53096 -11173 53247 -10830 0 FreeSans 480 270 0 0 VIN
port 26 nsew
flabel metal3 53497 -35185 53696 -34986 0 FreeSans 320 90 0 0 VCM
port 28 nsew
<< end >>
