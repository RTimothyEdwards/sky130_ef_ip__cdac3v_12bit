magic
tech sky130A
magscale 1 2
timestamp 1718225130
<< metal3 >>
rect 81341 -31712 81401 -31572
rect 81031 -32022 82511 -31712
rect 81031 -32082 82651 -32022
rect 81031 -32822 82511 -32082
rect 80891 -32882 82511 -32822
rect 81031 -33192 82511 -32882
rect 82141 -33332 82201 -33192
<< mimcap >>
rect 81071 -31792 82471 -31752
rect 81071 -33112 81111 -31792
rect 82431 -33112 82471 -31792
rect 81071 -33152 82471 -33112
<< mimcapcontact >>
rect 81111 -33112 82431 -31792
<< metal4 >>
rect 81741 -31672 81801 -31572
rect 80991 -31792 82551 -31672
rect 80991 -32422 81111 -31792
rect 80891 -32482 81111 -32422
rect 80991 -33112 81111 -32482
rect 82431 -32422 82551 -31792
rect 82431 -32482 82651 -32422
rect 82431 -33112 82551 -32482
rect 80991 -33232 82551 -33112
rect 81741 -33332 81801 -33232
<< mimcap2 >>
rect 81071 -31792 82471 -31752
rect 81071 -33112 81111 -31792
rect 82431 -33112 82471 -31792
rect 81071 -33152 82471 -33112
<< mimcap2contact >>
rect 81111 -33112 82431 -31792
<< metal5 >>
rect 82011 -31768 82331 -31077
rect 81087 -31792 82455 -31768
rect 81087 -31892 81111 -31792
rect 80396 -32212 81111 -31892
rect 81087 -33112 81111 -32212
rect 82431 -32692 82455 -31792
rect 82431 -33012 83146 -32692
rect 82431 -33112 82455 -33012
rect 81087 -33136 82455 -33112
rect 81211 -33828 81531 -33136
<< end >>
