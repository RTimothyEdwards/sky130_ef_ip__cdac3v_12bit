magic
tech sky130A
magscale 1 2
timestamp 1718247631
<< metal3 >>
rect 81341 -31713 81401 -31573
rect 81031 -32023 82511 -31713
rect 81031 -32083 82651 -32023
rect 81031 -32845 82511 -32083
rect 80891 -32905 82511 -32845
rect 81031 -33215 82511 -32905
rect 82141 -33355 82201 -33215
<< mimcap >>
rect 81071 -31793 82471 -31753
rect 81071 -33135 81111 -31793
rect 82431 -33135 82471 -31793
rect 81071 -33175 82471 -33135
<< mimcapcontact >>
rect 81111 -33135 82431 -31793
<< metal4 >>
rect 81741 -31673 81801 -31573
rect 80991 -31793 82551 -31673
rect 80991 -32434 81111 -31793
rect 80891 -32494 81111 -32434
rect 80991 -33135 81111 -32494
rect 82431 -32434 82551 -31793
rect 82431 -32494 82651 -32434
rect 82431 -33135 82551 -32494
rect 80991 -33255 82551 -33135
rect 81741 -33355 81801 -33255
<< mimcap2 >>
rect 81071 -31793 82471 -31753
rect 81071 -33135 81111 -31793
rect 82431 -33135 82471 -31793
rect 81071 -33175 82471 -33135
<< mimcap2contact >>
rect 81111 -33135 82431 -31793
<< metal5 >>
rect 82011 -31769 82331 -31078
rect 81087 -31793 82455 -31769
rect 81087 -31893 81111 -31793
rect 80396 -32213 81111 -31893
rect 81087 -33135 81111 -32213
rect 82431 -32715 82455 -31793
rect 82431 -33035 83146 -32715
rect 82431 -33135 82455 -33035
rect 81087 -33159 82455 -33135
rect 81211 -33851 81531 -33159
<< end >>
