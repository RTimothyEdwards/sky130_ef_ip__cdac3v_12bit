magic
tech sky130A
magscale 1 2
timestamp 1717891028
<< metal3 >>
rect -909 9172 909 9200
rect -909 7748 825 9172
rect 889 7748 909 9172
rect -909 7720 909 7748
rect -909 7372 909 7400
rect -909 5948 825 7372
rect 889 5948 909 7372
rect -909 5920 909 5948
rect -909 5572 909 5600
rect -909 4148 825 5572
rect 889 4148 909 5572
rect -909 4120 909 4148
rect -909 3772 909 3800
rect -909 2348 825 3772
rect 889 2348 909 3772
rect -909 2320 909 2348
rect -909 1972 909 2000
rect -909 548 825 1972
rect 889 548 909 1972
rect -909 520 909 548
rect -909 172 909 200
rect -909 -1252 825 172
rect 889 -1252 909 172
rect -909 -1280 909 -1252
rect -909 -1628 909 -1600
rect -909 -3052 825 -1628
rect 889 -3052 909 -1628
rect -909 -3080 909 -3052
rect -909 -3428 909 -3400
rect -909 -4852 825 -3428
rect 889 -4852 909 -3428
rect -909 -4880 909 -4852
rect -909 -5228 909 -5200
rect -909 -6652 825 -5228
rect 889 -6652 909 -5228
rect -909 -6680 909 -6652
rect -909 -7028 909 -7000
rect -909 -8452 825 -7028
rect 889 -8452 909 -7028
rect -909 -8480 909 -8452
<< via3 >>
rect 825 7748 889 9172
rect 825 5948 889 7372
rect 825 4148 889 5572
rect 825 2348 889 3772
rect 825 548 889 1972
rect 825 -1252 889 172
rect 825 -3052 889 -1628
rect 825 -4852 889 -3428
rect 825 -6652 889 -5228
rect 825 -8452 889 -7028
<< mimcap >>
rect -869 9120 577 9160
rect -869 7800 -829 9120
rect 537 7800 577 9120
rect -869 7760 577 7800
rect -869 7320 577 7360
rect -869 6000 -829 7320
rect 537 6000 577 7320
rect -869 5960 577 6000
rect -869 5520 577 5560
rect -869 4200 -829 5520
rect 537 4200 577 5520
rect -869 4160 577 4200
rect -869 3720 577 3760
rect -869 2400 -829 3720
rect 537 2400 577 3720
rect -869 2360 577 2400
rect -869 1920 577 1960
rect -869 600 -829 1920
rect 537 600 577 1920
rect -869 560 577 600
rect -869 120 577 160
rect -869 -1200 -829 120
rect 537 -1200 577 120
rect -869 -1240 577 -1200
rect -869 -1680 577 -1640
rect -869 -3000 -829 -1680
rect 537 -3000 577 -1680
rect -869 -3040 577 -3000
rect -869 -3480 577 -3440
rect -869 -4800 -829 -3480
rect 537 -4800 577 -3480
rect -869 -4840 577 -4800
rect -869 -5280 577 -5240
rect -869 -6600 -829 -5280
rect 537 -6600 577 -5280
rect -869 -6640 577 -6600
rect -869 -7080 577 -7040
rect -869 -8400 -829 -7080
rect 537 -8400 577 -7080
rect -869 -8440 577 -8400
<< mimcapcontact >>
rect -829 7800 537 9120
rect -829 6000 537 7320
rect -829 4200 537 5520
rect -829 2400 537 3720
rect -829 600 537 1920
rect -829 -1200 537 120
rect -829 -3000 537 -1680
rect -829 -4800 537 -3480
rect -829 -6600 537 -5280
rect -829 -8400 537 -7080
<< metal4 >>
rect 809 9172 905 9188
rect -830 9120 538 9121
rect -830 7800 -829 9120
rect 537 7800 538 9120
rect -830 7799 538 7800
rect 809 7748 825 9172
rect 889 7748 905 9172
rect 809 7732 905 7748
rect 809 7372 905 7388
rect -830 7320 538 7321
rect -830 6000 -829 7320
rect 537 6000 538 7320
rect -830 5999 538 6000
rect 809 5948 825 7372
rect 889 5948 905 7372
rect 809 5932 905 5948
rect 809 5572 905 5588
rect -830 5520 538 5521
rect -830 4200 -829 5520
rect 537 4200 538 5520
rect -830 4199 538 4200
rect 809 4148 825 5572
rect 889 4148 905 5572
rect 809 4132 905 4148
rect 809 3772 905 3788
rect -830 3720 538 3721
rect -830 2400 -829 3720
rect 537 2400 538 3720
rect -830 2399 538 2400
rect 809 2348 825 3772
rect 889 2348 905 3772
rect 809 2332 905 2348
rect 809 1972 905 1988
rect -830 1920 538 1921
rect -830 600 -829 1920
rect 537 600 538 1920
rect -830 599 538 600
rect 809 548 825 1972
rect 889 548 905 1972
rect 809 532 905 548
rect 809 172 905 188
rect -830 120 538 121
rect -830 -1200 -829 120
rect 537 -1200 538 120
rect -830 -1201 538 -1200
rect 809 -1252 825 172
rect 889 -1252 905 172
rect 809 -1268 905 -1252
rect 809 -1628 905 -1612
rect -830 -1680 538 -1679
rect -830 -3000 -829 -1680
rect 537 -3000 538 -1680
rect -830 -3001 538 -3000
rect 809 -3052 825 -1628
rect 889 -3052 905 -1628
rect 809 -3068 905 -3052
rect 809 -3428 905 -3412
rect -830 -3480 538 -3479
rect -830 -4800 -829 -3480
rect 537 -4800 538 -3480
rect -830 -4801 538 -4800
rect 809 -4852 825 -3428
rect 889 -4852 905 -3428
rect 809 -4868 905 -4852
rect 809 -5228 905 -5212
rect -830 -5280 538 -5279
rect -830 -6600 -829 -5280
rect 537 -6600 538 -5280
rect -830 -6601 538 -6600
rect 809 -6652 825 -5228
rect 889 -6652 905 -5228
rect 809 -6668 905 -6652
rect 809 -7028 905 -7012
rect -830 -7080 538 -7079
rect -830 -8400 -829 -7080
rect 537 -8400 538 -7080
rect -830 -8401 538 -8400
rect 809 -8452 825 -7028
rect 889 -8452 905 -7028
rect 809 -8468 905 -8452
<< properties >>
string FIXED_BBOX -909 7000 617 8480
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7.225 l 7.0 val 106.555 carea 2.00 cperi 0.19 nx 1 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
