magic
tech sky130A
magscale 1 2
timestamp 1718131540
<< locali >>
rect 3410 -3153 3810 -3137
rect 3410 -3324 3428 -3153
rect 3789 -3324 3810 -3153
rect 3410 -3340 3810 -3324
rect 4444 -5458 4557 -5457
rect 4556 -5492 4557 -5458
rect 4444 -5494 4557 -5492
rect 3409 -6990 3810 -6974
rect 3409 -7177 3426 -6990
rect 3794 -7177 3810 -6990
rect 3409 -7196 3810 -7177
<< viali >>
rect 3428 -3324 3789 -3153
rect 4444 -5492 4556 -5458
rect 4610 -5548 4644 -5412
rect 3426 -7177 3794 -6990
<< metal1 >>
rect 4880 -2560 5080 -2360
rect 3410 -3153 3810 -3137
rect 3410 -3324 3428 -3153
rect 3789 -3324 3810 -3153
rect 3410 -3340 3810 -3324
rect 4351 -3514 4551 -3513
rect 4126 -3662 4551 -3514
rect 4351 -3713 4551 -3662
rect 1240 -3925 3016 -3889
rect 656 -4196 856 -3996
rect 2980 -4009 3016 -3925
rect 4595 -4009 4601 -4001
rect 2980 -4045 4601 -4009
rect 4595 -4173 4601 -4045
rect 4653 -4173 4659 -4001
rect 673 -5265 873 -5065
rect 4113 -5290 4852 -5177
rect 4327 -5621 4333 -5447
rect 4385 -5458 4568 -5447
rect 4385 -5492 4444 -5458
rect 4556 -5492 4568 -5458
rect 4385 -5500 4568 -5492
rect 4385 -5621 4391 -5500
rect 4597 -5562 4603 -5390
rect 4655 -5562 4661 -5390
rect 666 -6104 1155 -5854
rect 4488 -6132 4603 -5738
rect 3195 -6189 4603 -6132
rect 4207 -6306 4213 -6298
rect 2901 -6342 4213 -6306
rect 2901 -6405 2937 -6342
rect 4207 -6350 4213 -6342
rect 4385 -6350 4391 -6298
rect 1224 -6441 2937 -6405
rect 666 -6729 866 -6529
rect 3409 -6990 3810 -6974
rect 3409 -7177 3426 -6990
rect 3794 -7177 3810 -6990
rect 3409 -7196 3810 -7177
rect 4880 -7970 5080 -7770
<< via1 >>
rect 2222 -1952 2596 -1833
rect 1628 -2855 1997 -2735
rect 3428 -3324 3789 -3153
rect 2098 -4198 2315 -4141
rect 2824 -4198 3201 -4141
rect 4601 -4173 4653 -4001
rect 3425 -5277 3795 -5051
rect 4333 -5621 4385 -5447
rect 4603 -5412 4655 -5390
rect 4603 -5548 4610 -5412
rect 4610 -5548 4644 -5412
rect 4644 -5548 4655 -5412
rect 4603 -5562 4655 -5548
rect 2098 -6189 2315 -6132
rect 2822 -6189 3195 -6132
rect 4213 -6350 4385 -6298
rect 3426 -7177 3794 -6990
rect 1622 -7598 1995 -7474
rect 2222 -8497 2597 -8374
<< metal2 >>
rect 2209 -1726 2610 -1712
rect 2209 -1952 2222 -1726
rect 2596 -1952 2610 -1726
rect 2209 -1965 2610 -1952
rect 1609 -2734 2010 -2722
rect 1609 -2945 1627 -2734
rect 1997 -2945 2010 -2734
rect 1609 -2956 2010 -2945
rect 3410 -3153 3810 -3137
rect 3410 -3324 3428 -3153
rect 3789 -3324 3810 -3153
rect 3410 -3340 3810 -3324
rect 4601 -4001 4653 -3995
rect 2812 -4063 3210 -4049
rect 2098 -4141 2315 -4132
rect 2812 -4198 2824 -4063
rect 3198 -4141 3210 -4063
rect 3201 -4198 3210 -4141
rect 4601 -4179 4653 -4173
rect 1279 -5859 1501 -4471
rect 2098 -6132 2315 -4198
rect 2468 -5860 2691 -4472
rect 3410 -5051 3809 -5040
rect 3410 -5277 3425 -5051
rect 3795 -5277 3809 -5051
rect 3410 -5290 3809 -5277
rect 4609 -5384 4645 -4179
rect 4603 -5390 4655 -5384
rect 4333 -5447 4385 -5441
rect 4603 -5568 4655 -5562
rect 4609 -5606 4645 -5568
rect 4333 -5627 4385 -5621
rect 2098 -6195 2315 -6189
rect 2810 -6148 2822 -6132
rect 2810 -6266 2821 -6148
rect 3195 -6266 3210 -6132
rect 2810 -6278 3210 -6266
rect 4341 -6292 4377 -5627
rect 4213 -6298 4385 -6292
rect 4213 -6356 4385 -6350
rect 3409 -6990 3810 -6974
rect 3409 -7177 3426 -6990
rect 3794 -7177 3810 -6990
rect 3409 -7196 3810 -7177
rect 1608 -7384 2010 -7369
rect 1608 -7598 1622 -7384
rect 1996 -7598 2010 -7384
rect 1608 -7607 2010 -7598
rect 2210 -8374 2610 -8364
rect 2210 -8375 2222 -8374
rect 2210 -8578 2221 -8375
rect 2597 -8578 2610 -8374
rect 2210 -8591 2610 -8578
<< via2 >>
rect 2222 -1833 2596 -1726
rect 2222 -1952 2596 -1833
rect 4600 -2320 4777 -2125
rect 1627 -2735 1997 -2734
rect 1627 -2855 1628 -2735
rect 1628 -2855 1997 -2735
rect 1627 -2945 1997 -2855
rect 3428 -3324 3789 -3153
rect 2824 -4141 3198 -4063
rect 2824 -4186 3198 -4141
rect 3425 -5277 3795 -5051
rect 2821 -6189 2822 -6148
rect 2822 -6189 3195 -6148
rect 2821 -6266 3195 -6189
rect 3426 -7177 3794 -6990
rect 1622 -7474 1996 -7384
rect 1622 -7598 1995 -7474
rect 1995 -7598 1996 -7474
rect 4600 -8205 4777 -8010
rect 2221 -8497 2222 -8375
rect 2222 -8497 2597 -8375
rect 2221 -8578 2597 -8497
<< metal3 >>
rect 1610 -2734 2010 -1606
rect 1610 -2945 1627 -2734
rect 1997 -2945 2010 -2734
rect 1610 -7384 2010 -2945
rect 1610 -7598 1622 -7384
rect 1996 -7598 2010 -7384
rect 1610 -8707 2010 -7598
rect 2210 -1726 2610 -1606
rect 2210 -1952 2222 -1726
rect 2596 -1952 2610 -1726
rect 2210 -8375 2610 -1952
rect 2210 -8578 2221 -8375
rect 2597 -8578 2610 -8375
rect 2210 -8707 2610 -8578
rect 2810 -4063 3210 -1598
rect 2810 -4186 2824 -4063
rect 3198 -4186 3210 -4063
rect 2810 -6148 3210 -4186
rect 2810 -6266 2821 -6148
rect 3195 -6266 3210 -6148
rect 2810 -8700 3210 -6266
rect 3410 -3153 3810 -1598
rect 3410 -3324 3428 -3153
rect 3789 -3324 3810 -3153
rect 3410 -5051 3810 -3324
rect 3410 -5277 3425 -5051
rect 3795 -5277 3810 -5051
rect 3410 -6990 3810 -5277
rect 3410 -7177 3426 -6990
rect 3794 -7177 3810 -6990
rect 3410 -8700 3810 -7177
rect 4591 -2125 4787 -2058
rect 4591 -2320 4600 -2125
rect 4777 -2320 4787 -2125
rect 4591 -6461 4787 -2320
rect 4591 -6661 4791 -6461
rect 4591 -8010 4787 -6661
rect 4591 -8205 4600 -8010
rect 4777 -8205 4787 -8010
rect 4591 -8254 4787 -8205
use simple_analog_switch_ena1v8  simple_analog_switch_ena1v8_1 ../dependencies/sky130_ef_ip__analog_switches/mag
timestamp 1718126855
transform 1 0 664 0 1 -8770
box 0 0 4416 3648
use simple_analog_switch_ena1v8  simple_analog_switch_ena1v8_2
timestamp 1718126855
transform 1 0 664 0 -1 -1560
box 0 0 4416 3648
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 4489 0 -1 -5242
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1715205430
transform 1 0 4765 0 -1 -5242
box -38 -48 130 592
<< labels >>
flabel metal1 673 -5265 873 -5065 0 FreeSans 256 0 0 0 dvss
port 7 nsew
flabel metal1 4351 -3713 4551 -3513 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 656 -4196 856 -3996 0 FreeSans 256 0 0 0 vdd1p8
port 1 nsew
flabel metal1 666 -6729 866 -6529 0 FreeSans 256 0 0 0 sel
port 6 nsew
flabel metal1 666 -6079 866 -5879 0 FreeSans 256 0 0 0 vdd3p3
port 0 nsew
flabel metal1 4880 -2560 5080 -2360 0 FreeSans 256 0 0 0 b
port 5 nsew
flabel metal1 4880 -7970 5080 -7770 0 FreeSans 256 0 0 0 a
port 4 nsew
flabel metal3 4591 -6661 4791 -6461 0 FreeSans 256 0 0 0 vo
port 2 nsew
<< end >>
