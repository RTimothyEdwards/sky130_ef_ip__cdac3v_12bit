magic
tech sky130A
magscale 1 2
timestamp 1722438219
<< viali >>
rect 58720 12899 83690 12933
rect 58631 -34472 58665 12845
rect 83747 -34470 83781 12837
rect 58722 -34559 83692 -34525
<< metal1 >>
rect 53524 14365 68765 14413
rect 53335 14269 70877 14317
rect 71172 14269 89082 14317
rect 53239 14173 69361 14221
rect 69662 14173 89177 14221
rect 53142 14077 70117 14125
rect 70415 14077 89273 14125
rect 53046 13981 72767 14029
rect 76033 13981 89368 14029
rect 76033 13933 76081 13981
rect 52949 13885 68727 13933
rect 72328 13885 76081 13933
rect 76152 13885 89464 13933
rect 68679 13837 68727 13885
rect 52849 13789 68605 13837
rect 68679 13789 72007 13837
rect 68557 13645 68605 13789
rect 76152 13741 76200 13885
rect 71570 13693 76200 13741
rect 76267 13789 89562 13837
rect 68557 13597 73528 13645
rect 76267 13549 76315 13789
rect 73085 13501 76315 13549
rect 58611 12933 83801 12953
rect 58611 12899 58720 12933
rect 83690 12899 83801 12933
rect 58611 12879 83801 12899
rect 58611 12845 58685 12879
rect 52856 8734 53526 8782
rect 52952 1730 53526 1778
rect 53048 -5275 53526 -5227
rect 53089 -19283 53526 -19235
rect 53089 -26286 53526 -26238
rect 53089 -33290 53526 -33242
rect 58611 -34472 58631 12845
rect 58665 -34472 58685 12845
rect 58611 -34505 58685 -34472
rect 83727 12837 83801 12879
rect 83727 -34470 83747 12837
rect 83781 -34470 83801 12837
rect 88887 8733 89557 8781
rect 88887 1730 89469 1778
rect 88887 -5274 89372 -5226
rect 88887 -19282 89306 -19234
rect 88886 -26286 89322 -26238
rect 88887 -33290 89322 -33242
rect 83727 -34505 83801 -34470
rect 58611 -34525 83801 -34505
rect 58611 -34559 58722 -34525
rect 83692 -34559 83801 -34525
rect 58611 -34579 83801 -34559
rect 58611 -34690 58685 -34579
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -34948 58685 -34939
rect 83727 -34698 83801 -34579
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 83727 -34955 83801 -34947
<< via1 >>
rect 58619 -34939 58678 -34690
rect 83734 -34947 83793 -34698
<< metal2 >>
rect 53488 14421 53565 14432
rect 52859 8730 52907 13786
rect 52955 1725 53003 13940
rect 53051 -5279 53099 14037
rect 53147 -19329 53195 14131
rect 53243 -26299 53291 14225
rect 53339 -33302 53387 14325
rect 53488 14235 53498 14421
rect 53555 14235 53565 14421
rect 53488 14224 53565 14235
rect 67192 13923 68325 14589
rect 68837 14413 69037 14589
rect 68765 14365 69037 14413
rect 69217 14389 69417 14589
rect 69602 14390 69802 14590
rect 69980 14391 70180 14591
rect 70363 14391 70563 14591
rect 70742 14391 70942 14591
rect 69294 14158 69342 14389
rect 69674 14158 69722 14390
rect 70054 14067 70102 14391
rect 70434 14067 70482 14391
rect 70814 14259 70862 14391
rect 71124 14389 71324 14589
rect 71501 14391 71701 14591
rect 71886 14391 72086 14591
rect 72256 14391 72456 14591
rect 72639 14391 72839 14591
rect 71194 14259 71242 14389
rect 67192 13577 67221 13923
rect 68290 13577 68325 13923
rect 71574 13692 71622 14391
rect 71954 13788 72002 14391
rect 72334 13881 72382 14391
rect 72714 13975 72762 14391
rect 73014 14389 73214 14589
rect 73392 14391 73592 14591
rect 74028 14498 75160 14592
rect 67192 13552 68325 13577
rect 73094 13494 73142 14389
rect 73474 13588 73522 14391
rect 74028 14149 74053 14498
rect 75137 14149 75160 14498
rect 74028 14123 75160 14149
rect 57639 -9376 57703 -7904
rect 53490 -9387 53561 -9377
rect 53490 -9561 53498 -9387
rect 53555 -9561 53561 -9387
rect 53490 -9570 53561 -9561
rect 57639 -9667 57703 -9658
rect 57639 -11972 57703 -11963
rect 57639 -13571 57703 -12254
rect 89029 -33326 89077 14327
rect 89125 -26323 89173 14226
rect 89221 -19307 89269 14132
rect 89317 -5309 89365 14033
rect 89413 1725 89461 13938
rect 89509 8726 89557 13844
rect 58611 -34690 58685 -34682
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -36347 58685 -34939
rect 83727 -34698 83801 -34690
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 68751 -35760 70341 -35717
rect 68751 -36098 68783 -35760
rect 70303 -36098 70341 -35760
rect 58611 -36358 58735 -36347
rect 58611 -36734 58624 -36358
rect 58724 -36734 58735 -36358
rect 58611 -36741 58735 -36734
rect 58612 -36746 58735 -36741
rect 68751 -36856 70341 -36098
rect 72201 -36381 73791 -36342
rect 83727 -36347 83801 -34947
rect 72201 -36719 72237 -36381
rect 73757 -36719 73791 -36381
rect 72201 -36868 73791 -36719
rect 83672 -36359 83801 -36347
rect 83672 -36735 83686 -36359
rect 83789 -36735 83801 -36359
rect 83672 -36747 83801 -36735
<< via2 >>
rect 53498 14235 53555 14421
rect 67221 13577 68290 13923
rect 74053 14149 75137 14498
rect 53498 -9561 53555 -9387
rect 57639 -9658 57703 -9376
rect 57639 -12254 57703 -11972
rect 68783 -36098 70303 -35760
rect 58624 -36734 58724 -36358
rect 72237 -36719 73757 -36381
rect 83686 -36735 83789 -36359
<< metal3 >>
rect 53488 14421 53565 14432
rect 53488 14235 53498 14421
rect 53555 14235 53565 14421
rect 53488 14224 53565 14235
rect 53496 -9377 53556 14224
rect 65040 14202 65240 14402
rect 64616 13678 64816 13878
rect 57444 10306 57452 10370
rect 57681 10306 58425 10370
rect 84059 10182 85236 10246
rect 57196 7826 58405 7890
rect 57189 2742 58413 2806
rect 83551 2742 84399 2806
rect 84606 2742 84613 2806
rect 83933 262 85241 326
rect 57199 -4698 58320 -4634
rect 85203 -6990 85398 -6851
rect 83918 -7054 85398 -6990
rect 57634 -9376 57708 -9370
rect 53490 -9387 53561 -9377
rect 53490 -9561 53498 -9387
rect 53555 -9561 53561 -9387
rect 53490 -9570 53561 -9561
rect 57634 -9658 57639 -9376
rect 57703 -9594 57708 -9376
rect 88726 -9586 88955 -9580
rect 84666 -9594 84873 -9588
rect 57703 -9658 58900 -9594
rect 83980 -9658 84671 -9594
rect 84867 -9658 84873 -9594
rect 57634 -9663 57708 -9658
rect 84666 -9664 84873 -9658
rect 88726 -9661 88735 -9586
rect 88946 -9594 88955 -9586
rect 89380 -9594 89580 -9508
rect 88946 -9658 89580 -9594
rect 88946 -9661 88955 -9658
rect 88726 -9668 88955 -9661
rect 89380 -9708 89580 -9658
rect 57634 -11972 57708 -11967
rect 57634 -12254 57639 -11972
rect 57703 -12036 58919 -11972
rect 83840 -12036 84037 -11972
rect 57703 -12254 57708 -12036
rect 57634 -12260 57708 -12254
rect 57014 -14640 58370 -14576
rect 57014 -14663 57210 -14640
rect 83950 -16996 85256 -16932
rect 57162 -21956 58447 -21892
rect 54633 -24342 55033 -24324
rect 54633 -24464 54649 -24342
rect 55017 -24464 55033 -24342
rect 58042 -24368 58280 -24356
rect 58042 -24434 58054 -24368
rect 58266 -24372 58280 -24368
rect 58266 -24434 58410 -24372
rect 58042 -24436 58410 -24434
rect 83988 -24436 85241 -24372
rect 58042 -24450 58280 -24436
rect 54633 -24480 55033 -24464
rect 83963 -29520 85239 -29456
rect 57194 -31876 58330 -31812
rect 83980 -32000 84409 -31936
rect 84644 -32000 84651 -31936
rect 70647 -35210 70847 -35010
rect 71047 -35490 71247 -35290
rect 65838 -36033 66038 -35833
rect 65303 -36648 65503 -36448
<< via3 >>
rect 54639 10282 55027 10405
rect 57452 10306 57681 10370
rect 84399 2742 84606 2806
rect 87392 2709 87769 2840
rect 84671 -9658 84867 -9594
rect 88735 -9661 88946 -9586
rect 54649 -24464 55017 -24342
rect 58054 -24434 58266 -24368
rect 84409 -32000 84644 -31936
rect 87386 -32019 87774 -31915
<< metal4 >>
rect 54633 10405 55033 10406
rect 54633 10282 54639 10405
rect 55027 10370 55033 10405
rect 57451 10370 57682 10371
rect 55027 10306 57452 10370
rect 57681 10306 57682 10370
rect 55027 10282 55033 10306
rect 57451 10305 57682 10306
rect 54633 10281 55033 10282
rect 87380 2840 87780 2851
rect 84398 2806 84607 2807
rect 87380 2806 87392 2840
rect 84398 2742 84399 2806
rect 84606 2742 87392 2806
rect 84398 2741 84607 2742
rect 87380 2709 87392 2742
rect 87769 2709 87780 2840
rect 87380 2697 87780 2709
rect 88726 -9586 88955 -9580
rect 84666 -9594 84873 -9588
rect 88726 -9594 88735 -9586
rect 84666 -9658 84671 -9594
rect 84867 -9658 88735 -9594
rect 84666 -9664 84873 -9658
rect 88726 -9661 88735 -9658
rect 88946 -9661 88955 -9586
rect 88726 -9668 88955 -9661
rect 54631 -24342 55037 -24324
rect 54631 -24464 54649 -24342
rect 55017 -24374 55037 -24342
rect 58042 -24368 58280 -24356
rect 58042 -24374 58054 -24368
rect 55017 -24434 58054 -24374
rect 58266 -24434 58280 -24368
rect 55017 -24464 55037 -24434
rect 58042 -24450 58280 -24434
rect 54631 -24480 55037 -24464
rect 87380 -31915 87780 -31914
rect 84408 -31936 84645 -31935
rect 87380 -31936 87386 -31915
rect 84408 -32000 84409 -31936
rect 84644 -32000 87386 -31936
rect 84408 -32001 84645 -32000
rect 87380 -32019 87386 -32000
rect 87774 -32019 87780 -31915
rect 87380 -32020 87780 -32019
use cdac_dummy_switch  cdac_dummy_switch_1
timestamp 1718247631
transform -1 0 133337 0 1 6988
box 44011 -15952 48431 -14149
use cdac_dummy_switch  cdac_dummy_switch_2
timestamp 1718247631
transform -1 0 133337 0 -1 -28520
box 44011 -15952 48431 -14149
use cdac_via_3cut  cdac_via_3cut_0
timestamp 1718247631
transform 1 0 212 0 1 34864
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_1
timestamp 1718247631
transform 1 0 597 0 1 -156
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_2
timestamp 1718247631
transform 1 0 501 0 1 6844
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_3
timestamp 1718247631
transform 1 0 405 0 1 13803
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_4
timestamp 1718247631
transform 1 0 308 0 1 27859
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_5
timestamp 1718247631
transform 1 0 36481 0 1 13852
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_6
timestamp 1718247631
transform 1 0 116 0 1 41869
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_7
timestamp 1718247631
transform 1 0 36286 0 1 -156
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_8
timestamp 1718247631
transform 1 0 36382 0 1 6846
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_9
timestamp 1718247631
transform 1 0 36571 0 1 27862
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_10
timestamp 1718247631
transform 1 0 36767 0 1 41869
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_11
timestamp 1718247631
transform 1 0 36670 0 1 34866
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_12
timestamp 1718247631
transform 1 0 116 0 1 46924
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_13
timestamp 1718247631
transform 1 0 213 0 1 47021
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_14
timestamp 1718247631
transform 1 0 308 0 1 47117
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_15
timestamp 1718247631
transform 1 0 404 0 1 47213
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_16
timestamp 1718247631
transform 1 0 501 0 1 47308
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_17
timestamp 1718247631
transform 1 0 595 0 1 47403
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_18
timestamp 1718247631
transform 1 0 36768 0 1 46925
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_19
timestamp 1718247631
transform 1 0 36670 0 1 47019
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_20
timestamp 1718247631
transform 1 0 36574 0 1 47117
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_21
timestamp 1718247631
transform 1 0 36478 0 1 47212
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_22
timestamp 1718247631
transform 1 0 36381 0 1 47309
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_23
timestamp 1718247631
transform 1 0 36286 0 1 47405
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_24
timestamp 1718247631
transform 0 1 103797 -1 0 67058
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_25
timestamp 1718247631
transform 0 1 102275 -1 0 66961
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_26
timestamp 1718247631
transform 0 1 104329 -1 0 67057
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_27
timestamp 1718247631
transform 0 1 103040 -1 0 66865
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_28
timestamp 1718247631
transform 0 1 102807 -1 0 66959
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_29
timestamp 1718247631
transform 0 1 103566 -1 0 66867
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_30
timestamp 1718247631
transform 0 1 104707 -1 0 66480
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_31
timestamp 1718247631
transform 0 1 105697 -1 0 66770
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_32
timestamp 1718247631
transform 0 1 105466 -1 0 66677
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_33
timestamp 1718247631
transform 0 1 104940 -1 0 66579
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_34
timestamp 1718247631
transform 0 1 106228 -1 0 66291
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_35
timestamp 1718247631
transform 0 1 106453 -1 0 66386
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_36
timestamp 1718247631
transform 0 1 86645 -1 0 67155
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_37
timestamp 1718247631
transform 0 1 101701 -1 0 67154
box 52740 -33138 52792 -32927
use EF_SW_RST  x1
timestamp 1722438116
transform 1 0 52769 0 -1 -10037
box 318 -2876 4934 4338
use EF_AMUX0201_ARRAY1  x3
timestamp 1722437419
transform 0 1 62083 -1 0 14841
box 320 -9004 51588 27251
use EF_BANK_CAP_12  x4
timestamp 1722438219
transform 1 0 0 0 1 -8000
box 58243 -26645 84124 21019
<< labels >>
flabel metal3 64616 13678 64816 13878 0 FreeSans 256 90 0 0 DVSS
port 12 nsew
flabel metal3 71047 -35490 71247 -35290 0 FreeSans 256 90 0 0 VH
port 14 nsew
flabel metal3 70647 -35210 70847 -35010 0 FreeSans 256 90 0 0 VL
port 15 nsew
flabel metal3 65838 -36033 66038 -35833 0 FreeSans 256 90 0 0 VSS
port 13 nsew
flabel metal3 65303 -36648 65503 -36448 0 FreeSans 256 90 0 0 VDD
port 10 nsew
flabel metal3 65040 14202 65240 14402 0 FreeSans 256 90 0 0 DVDD
port 11 nsew
flabel metal3 89380 -9708 89580 -9508 0 FreeSans 480 0 0 0 OUT
port 16 nsew
flabel metal2 71501 14391 71701 14591 0 FreeSans 480 0 0 0 SELD6
port 6 nsew
flabel metal2 73392 14391 73592 14591 0 FreeSans 480 0 0 0 SELD11
port 21 nsew
flabel metal2 73014 14389 73214 14589 0 FreeSans 480 0 0 0 SELD10
port 19 nsew
flabel metal2 72639 14391 72839 14591 0 FreeSans 480 0 0 0 SELD9
port 9 nsew
flabel metal2 71886 14391 72086 14591 0 FreeSans 480 0 0 0 SELD7
port 7 nsew
flabel metal2 72256 14391 72456 14591 0 FreeSans 480 0 0 0 SELD8
port 8 nsew
flabel metal2 69980 14391 70180 14591 0 FreeSans 480 0 0 0 SELD2
port 2 nsew
flabel metal2 70363 14391 70563 14591 0 FreeSans 480 0 0 0 SELD3
port 3 nsew
flabel metal2 70742 14391 70942 14591 0 FreeSans 480 0 0 0 SELD4
port 4 nsew
flabel metal2 71124 14389 71324 14589 0 FreeSans 480 0 0 0 SELD5
port 5 nsew
flabel metal2 69602 14390 69802 14590 0 FreeSans 480 0 0 0 SELD1
port 24 nsew
flabel metal2 69217 14389 69417 14589 0 FreeSans 480 0 0 0 SELD0
port 23 nsew
flabel metal2 68837 14389 69037 14589 0 FreeSans 480 0 0 0 RST
port 17 nsew
flabel metal3 83840 -12036 84037 -11972 0 FreeSans 480 0 0 0 OUTNC
port 22 nsew
<< end >>
