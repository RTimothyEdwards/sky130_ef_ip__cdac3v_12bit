magic
tech sky130A
magscale 1 2
timestamp 1718247631
<< error_p >>
rect 81108 -26399 81428 -26353
rect 81951 -26363 82185 -25907
rect 81108 -26635 81150 -26399
rect 81871 -26443 82265 -26363
rect 81871 -26507 82551 -26443
rect 81871 -26587 82265 -26507
rect 81108 -26673 81428 -26635
rect 81908 -26679 81950 -26587
rect 81908 -26721 82228 -26679
<< dnwell >>
rect 81951 -26507 82185 -26443
<< metal3 >>
rect 82038 -26443 82098 -26177
rect 80427 -26507 81151 -26443
rect 81385 -26507 82098 -26443
rect 82179 -26507 82908 -26443
rect 80427 -26631 81951 -26567
rect 82185 -26631 82908 -26567
rect 81238 -26897 81298 -26631
<< via3 >>
rect 81151 -26507 81385 -26443
rect 81951 -26631 82185 -26567
<< metal4 >>
rect 81950 -26443 82186 -26442
<< via4 >>
rect 81150 -26443 81386 -26399
rect 81150 -26507 81151 -26443
rect 81151 -26507 81385 -26443
rect 81385 -26507 81386 -26443
rect 81150 -26635 81386 -26507
rect 81950 -26567 82186 -26443
rect 81950 -26631 81951 -26567
rect 81951 -26631 82185 -26567
rect 82185 -26631 82186 -26567
rect 81950 -26679 82186 -26631
<< metal5 >>
rect 81108 -26399 81428 -26354
rect 81108 -26635 81150 -26399
rect 81386 -26635 81428 -26399
rect 81108 -26673 81428 -26635
rect 81908 -26443 82228 -26402
rect 81908 -26679 81950 -26443
rect 82186 -26679 82228 -26443
rect 81908 -26721 82228 -26679
<< end >>
