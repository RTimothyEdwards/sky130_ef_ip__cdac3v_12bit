magic
tech sky130A
magscale 1 2
timestamp 1718225130
<< error_p >>
rect 66120 -2290 66440 -2266
rect 66120 -2562 66144 -2290
rect 66120 -2586 66440 -2562
rect 66070 -3090 66390 -3066
rect 66070 -3362 66094 -3090
rect 66070 -3386 66390 -3362
<< metal3 >>
rect 66036 -2394 66100 -2388
rect 65895 -2456 66036 -2396
rect 66036 -2464 66100 -2458
rect 66411 -3194 66475 -3188
rect 66475 -3256 66615 -3196
rect 66411 -3264 66475 -3258
<< via3 >>
rect 66036 -2458 66100 -2394
rect 66411 -3258 66475 -3194
<< metal4 >>
rect 66035 -2394 66144 -2393
rect 66035 -2458 66036 -2394
rect 66100 -2458 66144 -2394
rect 66035 -2460 66144 -2458
rect 66225 -3090 66285 -2562
rect 66366 -3194 66476 -3193
rect 66366 -3258 66411 -3194
rect 66475 -3258 66476 -3194
rect 66366 -3259 66476 -3258
<< via4 >>
rect 66144 -2562 66416 -2290
rect 66094 -3362 66366 -3090
<< metal5 >>
rect 66120 -2290 66440 -2266
rect 66120 -2562 66144 -2290
rect 66416 -2562 66440 -2290
rect 66120 -2586 66440 -2562
rect 66070 -3090 66390 -3066
rect 66070 -3362 66094 -3090
rect 66366 -3362 66390 -3090
rect 66070 -3386 66390 -3362
<< end >>
