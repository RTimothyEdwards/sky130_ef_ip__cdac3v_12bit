magic
tech sky130A
magscale 1 2
timestamp 1717881426
<< error_p >>
rect 774 7319 1094 7401
rect 774 6999 1094 7081
rect 774 5519 1094 5601
rect 774 5199 1094 5281
rect 774 3719 1094 3801
rect 774 3399 1094 3481
rect 774 1919 1094 2001
rect 774 1599 1094 1681
rect 774 119 1094 201
rect 774 -201 1094 -119
rect 774 -1681 1094 -1599
rect 774 -2001 1094 -1919
rect 774 -3481 1094 -3399
rect 774 -3801 1094 -3719
rect 774 -5281 1094 -5199
rect 774 -5601 1094 -5519
rect 774 -7081 1094 -6999
rect 774 -7401 1094 -7319
<< metal4 >>
rect -1072 8839 1072 8880
rect -1072 7361 816 8839
rect 1052 7361 1072 8839
rect -1072 7320 1072 7361
rect -1072 7039 1072 7080
rect -1072 5561 816 7039
rect 1052 5561 1072 7039
rect -1072 5520 1072 5561
rect -1072 5239 1072 5280
rect -1072 3761 816 5239
rect 1052 3761 1072 5239
rect -1072 3720 1072 3761
rect -1072 3439 1072 3480
rect -1072 1961 816 3439
rect 1052 1961 1072 3439
rect -1072 1920 1072 1961
rect -1072 1639 1072 1680
rect -1072 161 816 1639
rect 1052 161 1072 1639
rect -1072 120 1072 161
rect -1072 -161 1072 -120
rect -1072 -1639 816 -161
rect 1052 -1639 1072 -161
rect -1072 -1680 1072 -1639
rect -1072 -1961 1072 -1920
rect -1072 -3439 816 -1961
rect 1052 -3439 1072 -1961
rect -1072 -3480 1072 -3439
rect -1072 -3761 1072 -3720
rect -1072 -5239 816 -3761
rect 1052 -5239 1072 -3761
rect -1072 -5280 1072 -5239
rect -1072 -5561 1072 -5520
rect -1072 -7039 816 -5561
rect 1052 -7039 1072 -5561
rect -1072 -7080 1072 -7039
rect -1072 -7361 1072 -7320
rect -1072 -8839 816 -7361
rect 1052 -8839 1072 -7361
rect -1072 -8880 1072 -8839
<< via4 >>
rect 816 7361 1052 8839
rect 816 5561 1052 7039
rect 816 3761 1052 5239
rect 816 1961 1052 3439
rect 816 161 1052 1639
rect 816 -1639 1052 -161
rect 816 -3439 1052 -1961
rect 816 -5239 1052 -3761
rect 816 -7039 1052 -5561
rect 816 -8839 1052 -7361
<< mimcap2 >>
rect -992 8760 454 8800
rect -992 7440 -952 8760
rect 414 7440 454 8760
rect -992 7400 454 7440
rect -992 6960 454 7000
rect -992 5640 -952 6960
rect 414 5640 454 6960
rect -992 5600 454 5640
rect -992 5160 454 5200
rect -992 3840 -952 5160
rect 414 3840 454 5160
rect -992 3800 454 3840
rect -992 3360 454 3400
rect -992 2040 -952 3360
rect 414 2040 454 3360
rect -992 2000 454 2040
rect -992 1560 454 1600
rect -992 240 -952 1560
rect 414 240 454 1560
rect -992 200 454 240
rect -992 -240 454 -200
rect -992 -1560 -952 -240
rect 414 -1560 454 -240
rect -992 -1600 454 -1560
rect -992 -2040 454 -2000
rect -992 -3360 -952 -2040
rect 414 -3360 454 -2040
rect -992 -3400 454 -3360
rect -992 -3840 454 -3800
rect -992 -5160 -952 -3840
rect 414 -5160 454 -3840
rect -992 -5200 454 -5160
rect -992 -5640 454 -5600
rect -992 -6960 -952 -5640
rect 414 -6960 454 -5640
rect -992 -7000 454 -6960
rect -992 -7440 454 -7400
rect -992 -8760 -952 -7440
rect 414 -8760 454 -7440
rect -992 -8800 454 -8760
<< mimcap2contact >>
rect -952 7440 414 8760
rect -952 5640 414 6960
rect -952 3840 414 5160
rect -952 2040 414 3360
rect -952 240 414 1560
rect -952 -1560 414 -240
rect -952 -3360 414 -2040
rect -952 -5160 414 -3840
rect -952 -6960 414 -5640
rect -952 -8760 414 -7440
<< metal5 >>
rect 774 8839 1094 8881
rect -976 8760 438 8784
rect -976 7440 -952 8760
rect 414 7440 438 8760
rect -976 7416 438 7440
rect 774 7361 816 8839
rect 1052 7361 1094 8839
rect 774 7319 1094 7361
rect 774 7039 1094 7081
rect -976 6960 438 6984
rect -976 5640 -952 6960
rect 414 5640 438 6960
rect -976 5616 438 5640
rect 774 5561 816 7039
rect 1052 5561 1094 7039
rect 774 5519 1094 5561
rect 774 5239 1094 5281
rect -976 5160 438 5184
rect -976 3840 -952 5160
rect 414 3840 438 5160
rect -976 3816 438 3840
rect 774 3761 816 5239
rect 1052 3761 1094 5239
rect 774 3719 1094 3761
rect 774 3439 1094 3481
rect -976 3360 438 3384
rect -976 2040 -952 3360
rect 414 2040 438 3360
rect -976 2016 438 2040
rect 774 1961 816 3439
rect 1052 1961 1094 3439
rect 774 1919 1094 1961
rect 774 1639 1094 1681
rect -976 1560 438 1584
rect -976 240 -952 1560
rect 414 240 438 1560
rect -976 216 438 240
rect 774 161 816 1639
rect 1052 161 1094 1639
rect 774 119 1094 161
rect 774 -161 1094 -119
rect -976 -240 438 -216
rect -976 -1560 -952 -240
rect 414 -1560 438 -240
rect -976 -1584 438 -1560
rect 774 -1639 816 -161
rect 1052 -1639 1094 -161
rect 774 -1681 1094 -1639
rect 774 -1961 1094 -1919
rect -976 -2040 438 -2016
rect -976 -3360 -952 -2040
rect 414 -3360 438 -2040
rect -976 -3384 438 -3360
rect 774 -3439 816 -1961
rect 1052 -3439 1094 -1961
rect 774 -3481 1094 -3439
rect 774 -3761 1094 -3719
rect -976 -3840 438 -3816
rect -976 -5160 -952 -3840
rect 414 -5160 438 -3840
rect -976 -5184 438 -5160
rect 774 -5239 816 -3761
rect 1052 -5239 1094 -3761
rect 774 -5281 1094 -5239
rect 774 -5561 1094 -5519
rect -976 -5640 438 -5616
rect -976 -6960 -952 -5640
rect 414 -6960 438 -5640
rect -976 -6984 438 -6960
rect 774 -7039 816 -5561
rect 1052 -7039 1094 -5561
rect 774 -7081 1094 -7039
rect 774 -7361 1094 -7319
rect -976 -7440 438 -7416
rect -976 -8760 -952 -7440
rect 414 -8760 438 -7440
rect -976 -8784 438 -8760
rect 774 -8839 816 -7361
rect 1052 -8839 1094 -7361
rect 774 -8881 1094 -8839
<< properties >>
string FIXED_BBOX -1072 7320 534 8880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 7.225 l 7.0 val 106.555 carea 2.00 cperi 0.19 nx 1 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
