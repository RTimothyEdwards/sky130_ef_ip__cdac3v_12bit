magic
tech sky130A
magscale 1 2
timestamp 1731117925
<< dnwell >>
rect 673 603 4874 1007
<< nwell >>
rect 634 2450 4105 2916
rect 737 2444 872 2450
rect 563 712 4983 904
rect 633 -1477 4104 -834
<< metal1 >>
rect 820 2564 961 2568
rect 820 2512 828 2564
rect 953 2541 961 2564
rect 953 2512 3127 2541
rect 820 2508 3127 2512
rect 820 2505 960 2508
rect 736 2473 3032 2477
rect 736 2421 742 2473
rect 867 2444 3032 2473
rect 867 2421 874 2444
rect 3094 2424 3127 2508
rect 736 2414 874 2421
rect 1267 2347 1663 2362
rect 1267 2086 1291 2347
rect 1639 2086 1663 2347
rect 1267 2065 1663 2086
rect 1866 1293 2266 1309
rect 1866 1069 1888 1293
rect 2239 1069 2266 1293
rect 1866 1054 2266 1069
rect 818 872 966 882
rect 818 818 819 872
rect 960 869 966 872
rect 1821 869 2021 944
rect 960 825 3127 869
rect 960 818 966 825
rect 1821 824 2021 825
rect 818 810 966 818
rect 737 746 919 748
rect 737 745 1823 746
rect 2023 745 3032 746
rect 737 744 3032 745
rect 737 692 744 744
rect 911 702 3032 744
rect 911 692 919 702
rect 737 687 919 692
rect 1265 615 1662 627
rect 1823 622 2023 702
rect 3083 669 3127 825
rect 1265 341 1279 615
rect 1652 341 1662 615
rect 1265 327 1662 341
rect 1864 -443 2264 -424
rect 1864 -626 1885 -443
rect 2243 -626 2264 -443
rect 1864 -650 2264 -626
<< via1 >>
rect 828 2512 953 2564
rect 742 2421 867 2473
rect 1291 2086 1639 2347
rect 1888 1069 2239 1293
rect 819 818 960 872
rect 744 692 911 744
rect 1279 341 1652 615
rect 1885 -626 2243 -443
<< metal2 >>
rect 820 2564 960 2568
rect 820 2512 828 2564
rect 953 2512 960 2564
rect 820 2505 960 2512
rect 736 2473 874 2477
rect 736 2421 742 2473
rect 867 2421 874 2473
rect 736 2414 874 2421
rect 737 748 775 2414
rect 916 2356 954 2505
rect 818 2318 954 2356
rect 1267 2347 1663 2362
rect 818 882 856 2318
rect 1267 2086 1291 2347
rect 1639 2086 1663 2347
rect 1267 2065 1663 2086
rect 4245 1793 4441 1894
rect 4245 1738 4252 1793
rect 4676 1704 4876 1904
rect 1866 1293 2266 1309
rect 1866 1069 1888 1293
rect 2239 1069 2266 1293
rect 1866 1054 2266 1069
rect 818 872 966 882
rect 818 818 819 872
rect 960 818 966 872
rect 818 810 966 818
rect 737 744 919 748
rect 737 692 744 744
rect 911 692 919 744
rect 737 687 919 692
rect 1265 615 1662 627
rect 1265 341 1279 615
rect 1652 341 1662 615
rect 1265 327 1662 341
rect 4257 10 4429 11
rect 4678 -274 4878 -74
rect 1864 -443 2264 -424
rect 1864 -626 1885 -443
rect 2243 -626 2264 -443
rect 1864 -650 2264 -626
<< via2 >>
rect 1291 2086 1639 2347
rect 4257 1511 4429 1641
rect 1888 1069 2239 1293
rect 1279 341 1652 615
rect 4257 11 4429 141
rect 1885 -626 2243 -443
<< metal3 >>
rect 1264 2347 1662 4328
rect 1264 2086 1291 2347
rect 1639 2086 1662 2347
rect 1264 615 1662 2086
rect 1264 341 1279 615
rect 1652 341 1662 615
rect 1264 -2874 1662 341
rect 1864 1293 2262 4326
rect 1864 1069 1888 1293
rect 2239 1069 2262 1293
rect 1864 -443 2262 1069
rect 2464 -194 2862 4338
rect 1864 -626 1885 -443
rect 2243 -626 2262 -443
rect 1864 -1700 2262 -626
rect 1864 -2876 2262 -2130
rect 2464 -2864 2862 -412
rect 3064 -2858 3464 4334
rect 4245 1641 4441 2857
rect 4245 1511 4257 1641
rect 4429 1511 4441 1641
rect 4245 141 4441 1511
rect 4245 11 4257 141
rect 4429 11 4441 141
rect 4245 -1207 4441 11
use simple_analog_switch  simple_analog_switch_0 ../dependencies/sky130_ef_ip__analog_switches/mag
timestamp 1722435879
transform 1 0 -14 0 1 -858
box 577 24 4997 1570
use simple_analog_switch  simple_analog_switch_1
timestamp 1722435879
transform 1 0 -14 0 1 880
box 577 24 4997 1570
<< labels >>
flabel metal3 3105 -1078 3305 -878 0 FreeSans 256 0 0 0 DVSS
port 6 nsew
flabel metal3 2539 -1067 2739 -867 0 FreeSans 256 0 0 0 DVDD
port 3 nsew
flabel metal3 1938 -1037 2138 -891 0 FreeSans 256 0 0 0 AVSS
port 4 nsew
flabel metal3 1375 -1043 1575 -843 0 FreeSans 256 0 0 0 AVDD
port 2 nsew
flabel metal3 4245 712 4441 904 0 FreeSans 480 0 0 0 VIN
port 11 nsew
flabel metal2 4676 1704 4876 1904 0 FreeSans 256 0 0 0 VP1
port 1 nsew
flabel metal2 4678 -274 4878 -74 0 FreeSans 256 0 0 0 VP2
port 0 nsew
flabel metal1 1821 824 2021 944 0 FreeSans 256 0 0 0 HOLD
port 5 nsew
flabel metal1 1823 622 2023 745 0 FreeSans 320 0 0 0 HOLDB
port 10 nsew
<< end >>
