magic
tech sky130A
magscale 1 2
timestamp 1717890828
<< metal3 >>
rect -8934 9172 -7162 9200
rect -8934 7748 -7246 9172
rect -7182 7748 -7162 9172
rect -8934 7720 -7162 7748
rect -6436 9172 -4664 9200
rect -6436 7748 -4748 9172
rect -4684 7748 -4664 9172
rect -6436 7720 -4664 7748
rect -3938 9172 -2166 9200
rect -3938 7748 -2250 9172
rect -2186 7748 -2166 9172
rect -3938 7720 -2166 7748
rect -1440 9172 332 9200
rect -1440 7748 248 9172
rect 312 7748 332 9172
rect -1440 7720 332 7748
rect 1058 9172 2830 9200
rect 1058 7748 2746 9172
rect 2810 7748 2830 9172
rect 1058 7720 2830 7748
rect 3556 9172 5328 9200
rect 3556 7748 5244 9172
rect 5308 7748 5328 9172
rect 3556 7720 5328 7748
rect 6054 9172 7826 9200
rect 6054 7748 7742 9172
rect 7806 7748 7826 9172
rect 6054 7720 7826 7748
rect 8552 9172 10324 9200
rect 8552 7748 10240 9172
rect 10304 7748 10324 9172
rect 8552 7720 10324 7748
rect 11050 9172 12822 9200
rect 11050 7748 12738 9172
rect 12802 7748 12822 9172
rect 11050 7720 12822 7748
rect -8934 7372 -7162 7400
rect -8934 5948 -7246 7372
rect -7182 5948 -7162 7372
rect -8934 5920 -7162 5948
rect -6436 7372 -4664 7400
rect -6436 5948 -4748 7372
rect -4684 5948 -4664 7372
rect -6436 5920 -4664 5948
rect -3938 7372 -2166 7400
rect -3938 5948 -2250 7372
rect -2186 5948 -2166 7372
rect -3938 5920 -2166 5948
rect -1440 7372 332 7400
rect -1440 5948 248 7372
rect 312 5948 332 7372
rect -1440 5920 332 5948
rect 1058 7372 2830 7400
rect 1058 5948 2746 7372
rect 2810 5948 2830 7372
rect 1058 5920 2830 5948
rect 3556 7372 5328 7400
rect 3556 5948 5244 7372
rect 5308 5948 5328 7372
rect 3556 5920 5328 5948
rect 6054 7372 7826 7400
rect 6054 5948 7742 7372
rect 7806 5948 7826 7372
rect 6054 5920 7826 5948
rect 8552 7372 10324 7400
rect 8552 5948 10240 7372
rect 10304 5948 10324 7372
rect 8552 5920 10324 5948
rect 11050 7372 12822 7400
rect 11050 5948 12738 7372
rect 12802 5948 12822 7372
rect 11050 5920 12822 5948
rect -8934 5572 -7162 5600
rect -8934 4148 -7246 5572
rect -7182 4148 -7162 5572
rect -8934 4120 -7162 4148
rect -6436 5572 -4664 5600
rect -6436 4148 -4748 5572
rect -4684 4148 -4664 5572
rect -6436 4120 -4664 4148
rect -3938 5572 -2166 5600
rect -3938 4148 -2250 5572
rect -2186 4148 -2166 5572
rect -3938 4120 -2166 4148
rect -1440 5572 332 5600
rect -1440 4148 248 5572
rect 312 4148 332 5572
rect -1440 4120 332 4148
rect 1058 5572 2830 5600
rect 1058 4148 2746 5572
rect 2810 4148 2830 5572
rect 1058 4120 2830 4148
rect 3556 5572 5328 5600
rect 3556 4148 5244 5572
rect 5308 4148 5328 5572
rect 3556 4120 5328 4148
rect 6054 5572 7826 5600
rect 6054 4148 7742 5572
rect 7806 4148 7826 5572
rect 6054 4120 7826 4148
rect 8552 5572 10324 5600
rect 8552 4148 10240 5572
rect 10304 4148 10324 5572
rect 8552 4120 10324 4148
rect 11050 5572 12822 5600
rect 11050 4148 12738 5572
rect 12802 4148 12822 5572
rect 11050 4120 12822 4148
rect -8934 3772 -7162 3800
rect -8934 2348 -7246 3772
rect -7182 2348 -7162 3772
rect -8934 2320 -7162 2348
rect -6436 3772 -4664 3800
rect -6436 2348 -4748 3772
rect -4684 2348 -4664 3772
rect -6436 2320 -4664 2348
rect -3938 3772 -2166 3800
rect -3938 2348 -2250 3772
rect -2186 2348 -2166 3772
rect -3938 2320 -2166 2348
rect -1440 3772 332 3800
rect -1440 2348 248 3772
rect 312 2348 332 3772
rect -1440 2320 332 2348
rect 1058 3772 2830 3800
rect 1058 2348 2746 3772
rect 2810 2348 2830 3772
rect 1058 2320 2830 2348
rect 3556 3772 5328 3800
rect 3556 2348 5244 3772
rect 5308 2348 5328 3772
rect 3556 2320 5328 2348
rect 6054 3772 7826 3800
rect 6054 2348 7742 3772
rect 7806 2348 7826 3772
rect 6054 2320 7826 2348
rect 8552 3772 10324 3800
rect 8552 2348 10240 3772
rect 10304 2348 10324 3772
rect 8552 2320 10324 2348
rect 11050 3772 12822 3800
rect 11050 2348 12738 3772
rect 12802 2348 12822 3772
rect 11050 2320 12822 2348
rect -8934 1972 -7162 2000
rect -8934 548 -7246 1972
rect -7182 548 -7162 1972
rect -8934 520 -7162 548
rect -6436 1972 -4664 2000
rect -6436 548 -4748 1972
rect -4684 548 -4664 1972
rect -6436 520 -4664 548
rect -3938 1972 -2166 2000
rect -3938 548 -2250 1972
rect -2186 548 -2166 1972
rect -3938 520 -2166 548
rect -1440 1972 332 2000
rect -1440 548 248 1972
rect 312 548 332 1972
rect -1440 520 332 548
rect 1058 1972 2830 2000
rect 1058 548 2746 1972
rect 2810 548 2830 1972
rect 1058 520 2830 548
rect 3556 1972 5328 2000
rect 3556 548 5244 1972
rect 5308 548 5328 1972
rect 3556 520 5328 548
rect 6054 1972 7826 2000
rect 6054 548 7742 1972
rect 7806 548 7826 1972
rect 6054 520 7826 548
rect 8552 1972 10324 2000
rect 8552 548 10240 1972
rect 10304 548 10324 1972
rect 8552 520 10324 548
rect 11050 1972 12822 2000
rect 11050 548 12738 1972
rect 12802 548 12822 1972
rect 11050 520 12822 548
rect -8934 172 -7162 200
rect -8934 -1252 -7246 172
rect -7182 -1252 -7162 172
rect -8934 -1280 -7162 -1252
rect -6436 172 -4664 200
rect -6436 -1252 -4748 172
rect -4684 -1252 -4664 172
rect -6436 -1280 -4664 -1252
rect -3938 172 -2166 200
rect -3938 -1252 -2250 172
rect -2186 -1252 -2166 172
rect -3938 -1280 -2166 -1252
rect -1440 172 332 200
rect -1440 -1252 248 172
rect 312 -1252 332 172
rect -1440 -1280 332 -1252
rect 1058 172 2830 200
rect 1058 -1252 2746 172
rect 2810 -1252 2830 172
rect 1058 -1280 2830 -1252
rect 3556 172 5328 200
rect 3556 -1252 5244 172
rect 5308 -1252 5328 172
rect 3556 -1280 5328 -1252
rect 6054 172 7826 200
rect 6054 -1252 7742 172
rect 7806 -1252 7826 172
rect 6054 -1280 7826 -1252
rect 8552 172 10324 200
rect 8552 -1252 10240 172
rect 10304 -1252 10324 172
rect 8552 -1280 10324 -1252
rect 11050 172 12822 200
rect 11050 -1252 12738 172
rect 12802 -1252 12822 172
rect 11050 -1280 12822 -1252
rect -8934 -1628 -7162 -1600
rect -8934 -3052 -7246 -1628
rect -7182 -3052 -7162 -1628
rect -8934 -3080 -7162 -3052
rect -6436 -1628 -4664 -1600
rect -6436 -3052 -4748 -1628
rect -4684 -3052 -4664 -1628
rect -6436 -3080 -4664 -3052
rect -3938 -1628 -2166 -1600
rect -3938 -3052 -2250 -1628
rect -2186 -3052 -2166 -1628
rect -3938 -3080 -2166 -3052
rect -1440 -1628 332 -1600
rect -1440 -3052 248 -1628
rect 312 -3052 332 -1628
rect -1440 -3080 332 -3052
rect 1058 -1628 2830 -1600
rect 1058 -3052 2746 -1628
rect 2810 -3052 2830 -1628
rect 1058 -3080 2830 -3052
rect 3556 -1628 5328 -1600
rect 3556 -3052 5244 -1628
rect 5308 -3052 5328 -1628
rect 3556 -3080 5328 -3052
rect 6054 -1628 7826 -1600
rect 6054 -3052 7742 -1628
rect 7806 -3052 7826 -1628
rect 6054 -3080 7826 -3052
rect 8552 -1628 10324 -1600
rect 8552 -3052 10240 -1628
rect 10304 -3052 10324 -1628
rect 8552 -3080 10324 -3052
rect 11050 -1628 12822 -1600
rect 11050 -3052 12738 -1628
rect 12802 -3052 12822 -1628
rect 11050 -3080 12822 -3052
rect -8934 -3428 -7162 -3400
rect -8934 -4852 -7246 -3428
rect -7182 -4852 -7162 -3428
rect -8934 -4880 -7162 -4852
rect -6436 -3428 -4664 -3400
rect -6436 -4852 -4748 -3428
rect -4684 -4852 -4664 -3428
rect -6436 -4880 -4664 -4852
rect -3938 -3428 -2166 -3400
rect -3938 -4852 -2250 -3428
rect -2186 -4852 -2166 -3428
rect -3938 -4880 -2166 -4852
rect -1440 -3428 332 -3400
rect -1440 -4852 248 -3428
rect 312 -4852 332 -3428
rect -1440 -4880 332 -4852
rect 1058 -3428 2830 -3400
rect 1058 -4852 2746 -3428
rect 2810 -4852 2830 -3428
rect 1058 -4880 2830 -4852
rect 3556 -3428 5328 -3400
rect 3556 -4852 5244 -3428
rect 5308 -4852 5328 -3428
rect 3556 -4880 5328 -4852
rect 6054 -3428 7826 -3400
rect 6054 -4852 7742 -3428
rect 7806 -4852 7826 -3428
rect 6054 -4880 7826 -4852
rect 8552 -3428 10324 -3400
rect 8552 -4852 10240 -3428
rect 10304 -4852 10324 -3428
rect 8552 -4880 10324 -4852
rect 11050 -3428 12822 -3400
rect 11050 -4852 12738 -3428
rect 12802 -4852 12822 -3428
rect 11050 -4880 12822 -4852
rect -8934 -5228 -7162 -5200
rect -8934 -6652 -7246 -5228
rect -7182 -6652 -7162 -5228
rect -8934 -6680 -7162 -6652
rect -6436 -5228 -4664 -5200
rect -6436 -6652 -4748 -5228
rect -4684 -6652 -4664 -5228
rect -6436 -6680 -4664 -6652
rect -3938 -5228 -2166 -5200
rect -3938 -6652 -2250 -5228
rect -2186 -6652 -2166 -5228
rect -3938 -6680 -2166 -6652
rect -1440 -5228 332 -5200
rect -1440 -6652 248 -5228
rect 312 -6652 332 -5228
rect -1440 -6680 332 -6652
rect 1058 -5228 2830 -5200
rect 1058 -6652 2746 -5228
rect 2810 -6652 2830 -5228
rect 1058 -6680 2830 -6652
rect 3556 -5228 5328 -5200
rect 3556 -6652 5244 -5228
rect 5308 -6652 5328 -5228
rect 3556 -6680 5328 -6652
rect 6054 -5228 7826 -5200
rect 6054 -6652 7742 -5228
rect 7806 -6652 7826 -5228
rect 6054 -6680 7826 -6652
rect 8552 -5228 10324 -5200
rect 8552 -6652 10240 -5228
rect 10304 -6652 10324 -5228
rect 8552 -6680 10324 -6652
rect 11050 -5228 12822 -5200
rect 11050 -6652 12738 -5228
rect 12802 -6652 12822 -5228
rect 11050 -6680 12822 -6652
rect -8934 -7028 -7162 -7000
rect -8934 -8452 -7246 -7028
rect -7182 -8452 -7162 -7028
rect -8934 -8480 -7162 -8452
rect -6436 -7028 -4664 -7000
rect -6436 -8452 -4748 -7028
rect -4684 -8452 -4664 -7028
rect -6436 -8480 -4664 -8452
rect -3938 -7028 -2166 -7000
rect -3938 -8452 -2250 -7028
rect -2186 -8452 -2166 -7028
rect -3938 -8480 -2166 -8452
rect -1440 -7028 332 -7000
rect -1440 -8452 248 -7028
rect 312 -8452 332 -7028
rect -1440 -8480 332 -8452
rect 1058 -7028 2830 -7000
rect 1058 -8452 2746 -7028
rect 2810 -8452 2830 -7028
rect 1058 -8480 2830 -8452
rect 3556 -7028 5328 -7000
rect 3556 -8452 5244 -7028
rect 5308 -8452 5328 -7028
rect 3556 -8480 5328 -8452
rect 6054 -7028 7826 -7000
rect 6054 -8452 7742 -7028
rect 7806 -8452 7826 -7028
rect 6054 -8480 7826 -8452
rect 8552 -7028 10324 -7000
rect 8552 -8452 10240 -7028
rect 10304 -8452 10324 -7028
rect 8552 -8480 10324 -8452
rect 11050 -7028 12822 -7000
rect 11050 -8452 12738 -7028
rect 12802 -8452 12822 -7028
rect 11050 -8480 12822 -8452
<< via3 >>
rect -7246 7748 -7182 9172
rect -4748 7748 -4684 9172
rect -2250 7748 -2186 9172
rect 248 7748 312 9172
rect 2746 7748 2810 9172
rect 5244 7748 5308 9172
rect 7742 7748 7806 9172
rect 10240 7748 10304 9172
rect 12738 7748 12802 9172
rect -7246 5948 -7182 7372
rect -4748 5948 -4684 7372
rect -2250 5948 -2186 7372
rect 248 5948 312 7372
rect 2746 5948 2810 7372
rect 5244 5948 5308 7372
rect 7742 5948 7806 7372
rect 10240 5948 10304 7372
rect 12738 5948 12802 7372
rect -7246 4148 -7182 5572
rect -4748 4148 -4684 5572
rect -2250 4148 -2186 5572
rect 248 4148 312 5572
rect 2746 4148 2810 5572
rect 5244 4148 5308 5572
rect 7742 4148 7806 5572
rect 10240 4148 10304 5572
rect 12738 4148 12802 5572
rect -7246 2348 -7182 3772
rect -4748 2348 -4684 3772
rect -2250 2348 -2186 3772
rect 248 2348 312 3772
rect 2746 2348 2810 3772
rect 5244 2348 5308 3772
rect 7742 2348 7806 3772
rect 10240 2348 10304 3772
rect 12738 2348 12802 3772
rect -7246 548 -7182 1972
rect -4748 548 -4684 1972
rect -2250 548 -2186 1972
rect 248 548 312 1972
rect 2746 548 2810 1972
rect 5244 548 5308 1972
rect 7742 548 7806 1972
rect 10240 548 10304 1972
rect 12738 548 12802 1972
rect -7246 -1252 -7182 172
rect -4748 -1252 -4684 172
rect -2250 -1252 -2186 172
rect 248 -1252 312 172
rect 2746 -1252 2810 172
rect 5244 -1252 5308 172
rect 7742 -1252 7806 172
rect 10240 -1252 10304 172
rect 12738 -1252 12802 172
rect -7246 -3052 -7182 -1628
rect -4748 -3052 -4684 -1628
rect -2250 -3052 -2186 -1628
rect 248 -3052 312 -1628
rect 2746 -3052 2810 -1628
rect 5244 -3052 5308 -1628
rect 7742 -3052 7806 -1628
rect 10240 -3052 10304 -1628
rect 12738 -3052 12802 -1628
rect -7246 -4852 -7182 -3428
rect -4748 -4852 -4684 -3428
rect -2250 -4852 -2186 -3428
rect 248 -4852 312 -3428
rect 2746 -4852 2810 -3428
rect 5244 -4852 5308 -3428
rect 7742 -4852 7806 -3428
rect 10240 -4852 10304 -3428
rect 12738 -4852 12802 -3428
rect -7246 -6652 -7182 -5228
rect -4748 -6652 -4684 -5228
rect -2250 -6652 -2186 -5228
rect 248 -6652 312 -5228
rect 2746 -6652 2810 -5228
rect 5244 -6652 5308 -5228
rect 7742 -6652 7806 -5228
rect 10240 -6652 10304 -5228
rect 12738 -6652 12802 -5228
rect -7246 -8452 -7182 -7028
rect -4748 -8452 -4684 -7028
rect -2250 -8452 -2186 -7028
rect 248 -8452 312 -7028
rect 2746 -8452 2810 -7028
rect 5244 -8452 5308 -7028
rect 7742 -8452 7806 -7028
rect 10240 -8452 10304 -7028
rect 12738 -8452 12802 -7028
<< mimcap >>
rect -8894 9120 -7494 9160
rect -8894 7800 -8854 9120
rect -7534 7800 -7494 9120
rect -8894 7760 -7494 7800
rect -6396 9120 -4996 9160
rect -6396 7800 -6356 9120
rect -5036 7800 -4996 9120
rect -6396 7760 -4996 7800
rect -3898 9120 -2498 9160
rect -3898 7800 -3858 9120
rect -2538 7800 -2498 9120
rect -3898 7760 -2498 7800
rect -1400 9120 0 9160
rect -1400 7800 -1360 9120
rect -40 7800 0 9120
rect -1400 7760 0 7800
rect 1098 9120 2498 9160
rect 1098 7800 1138 9120
rect 2458 7800 2498 9120
rect 1098 7760 2498 7800
rect 3596 9120 4996 9160
rect 3596 7800 3636 9120
rect 4956 7800 4996 9120
rect 3596 7760 4996 7800
rect 6094 9120 7494 9160
rect 6094 7800 6134 9120
rect 7454 7800 7494 9120
rect 6094 7760 7494 7800
rect 8592 9120 9992 9160
rect 8592 7800 8632 9120
rect 9952 7800 9992 9120
rect 8592 7760 9992 7800
rect 11090 9120 12490 9160
rect 11090 7800 11130 9120
rect 12450 7800 12490 9120
rect 11090 7760 12490 7800
rect -8894 7320 -7494 7360
rect -8894 6000 -8854 7320
rect -7534 6000 -7494 7320
rect -8894 5960 -7494 6000
rect -6396 7320 -4996 7360
rect -6396 6000 -6356 7320
rect -5036 6000 -4996 7320
rect -6396 5960 -4996 6000
rect -3898 7320 -2498 7360
rect -3898 6000 -3858 7320
rect -2538 6000 -2498 7320
rect -3898 5960 -2498 6000
rect -1400 7320 0 7360
rect -1400 6000 -1360 7320
rect -40 6000 0 7320
rect -1400 5960 0 6000
rect 1098 7320 2498 7360
rect 1098 6000 1138 7320
rect 2458 6000 2498 7320
rect 1098 5960 2498 6000
rect 3596 7320 4996 7360
rect 3596 6000 3636 7320
rect 4956 6000 4996 7320
rect 3596 5960 4996 6000
rect 6094 7320 7494 7360
rect 6094 6000 6134 7320
rect 7454 6000 7494 7320
rect 6094 5960 7494 6000
rect 8592 7320 9992 7360
rect 8592 6000 8632 7320
rect 9952 6000 9992 7320
rect 8592 5960 9992 6000
rect 11090 7320 12490 7360
rect 11090 6000 11130 7320
rect 12450 6000 12490 7320
rect 11090 5960 12490 6000
rect -8894 5520 -7494 5560
rect -8894 4200 -8854 5520
rect -7534 4200 -7494 5520
rect -8894 4160 -7494 4200
rect -6396 5520 -4996 5560
rect -6396 4200 -6356 5520
rect -5036 4200 -4996 5520
rect -6396 4160 -4996 4200
rect -3898 5520 -2498 5560
rect -3898 4200 -3858 5520
rect -2538 4200 -2498 5520
rect -3898 4160 -2498 4200
rect -1400 5520 0 5560
rect -1400 4200 -1360 5520
rect -40 4200 0 5520
rect -1400 4160 0 4200
rect 1098 5520 2498 5560
rect 1098 4200 1138 5520
rect 2458 4200 2498 5520
rect 1098 4160 2498 4200
rect 3596 5520 4996 5560
rect 3596 4200 3636 5520
rect 4956 4200 4996 5520
rect 3596 4160 4996 4200
rect 6094 5520 7494 5560
rect 6094 4200 6134 5520
rect 7454 4200 7494 5520
rect 6094 4160 7494 4200
rect 8592 5520 9992 5560
rect 8592 4200 8632 5520
rect 9952 4200 9992 5520
rect 8592 4160 9992 4200
rect 11090 5520 12490 5560
rect 11090 4200 11130 5520
rect 12450 4200 12490 5520
rect 11090 4160 12490 4200
rect -8894 3720 -7494 3760
rect -8894 2400 -8854 3720
rect -7534 2400 -7494 3720
rect -8894 2360 -7494 2400
rect -6396 3720 -4996 3760
rect -6396 2400 -6356 3720
rect -5036 2400 -4996 3720
rect -6396 2360 -4996 2400
rect -3898 3720 -2498 3760
rect -3898 2400 -3858 3720
rect -2538 2400 -2498 3720
rect -3898 2360 -2498 2400
rect -1400 3720 0 3760
rect -1400 2400 -1360 3720
rect -40 2400 0 3720
rect -1400 2360 0 2400
rect 1098 3720 2498 3760
rect 1098 2400 1138 3720
rect 2458 2400 2498 3720
rect 1098 2360 2498 2400
rect 3596 3720 4996 3760
rect 3596 2400 3636 3720
rect 4956 2400 4996 3720
rect 3596 2360 4996 2400
rect 6094 3720 7494 3760
rect 6094 2400 6134 3720
rect 7454 2400 7494 3720
rect 6094 2360 7494 2400
rect 8592 3720 9992 3760
rect 8592 2400 8632 3720
rect 9952 2400 9992 3720
rect 8592 2360 9992 2400
rect 11090 3720 12490 3760
rect 11090 2400 11130 3720
rect 12450 2400 12490 3720
rect 11090 2360 12490 2400
rect -8894 1920 -7494 1960
rect -8894 600 -8854 1920
rect -7534 600 -7494 1920
rect -8894 560 -7494 600
rect -6396 1920 -4996 1960
rect -6396 600 -6356 1920
rect -5036 600 -4996 1920
rect -6396 560 -4996 600
rect -3898 1920 -2498 1960
rect -3898 600 -3858 1920
rect -2538 600 -2498 1920
rect -3898 560 -2498 600
rect -1400 1920 0 1960
rect -1400 600 -1360 1920
rect -40 600 0 1920
rect -1400 560 0 600
rect 1098 1920 2498 1960
rect 1098 600 1138 1920
rect 2458 600 2498 1920
rect 1098 560 2498 600
rect 3596 1920 4996 1960
rect 3596 600 3636 1920
rect 4956 600 4996 1920
rect 3596 560 4996 600
rect 6094 1920 7494 1960
rect 6094 600 6134 1920
rect 7454 600 7494 1920
rect 6094 560 7494 600
rect 8592 1920 9992 1960
rect 8592 600 8632 1920
rect 9952 600 9992 1920
rect 8592 560 9992 600
rect 11090 1920 12490 1960
rect 11090 600 11130 1920
rect 12450 600 12490 1920
rect 11090 560 12490 600
rect -8894 120 -7494 160
rect -8894 -1200 -8854 120
rect -7534 -1200 -7494 120
rect -8894 -1240 -7494 -1200
rect -6396 120 -4996 160
rect -6396 -1200 -6356 120
rect -5036 -1200 -4996 120
rect -6396 -1240 -4996 -1200
rect -3898 120 -2498 160
rect -3898 -1200 -3858 120
rect -2538 -1200 -2498 120
rect -3898 -1240 -2498 -1200
rect -1400 120 0 160
rect -1400 -1200 -1360 120
rect -40 -1200 0 120
rect -1400 -1240 0 -1200
rect 1098 120 2498 160
rect 1098 -1200 1138 120
rect 2458 -1200 2498 120
rect 1098 -1240 2498 -1200
rect 3596 120 4996 160
rect 3596 -1200 3636 120
rect 4956 -1200 4996 120
rect 3596 -1240 4996 -1200
rect 6094 120 7494 160
rect 6094 -1200 6134 120
rect 7454 -1200 7494 120
rect 6094 -1240 7494 -1200
rect 8592 120 9992 160
rect 8592 -1200 8632 120
rect 9952 -1200 9992 120
rect 8592 -1240 9992 -1200
rect 11090 120 12490 160
rect 11090 -1200 11130 120
rect 12450 -1200 12490 120
rect 11090 -1240 12490 -1200
rect -8894 -1680 -7494 -1640
rect -8894 -3000 -8854 -1680
rect -7534 -3000 -7494 -1680
rect -8894 -3040 -7494 -3000
rect -6396 -1680 -4996 -1640
rect -6396 -3000 -6356 -1680
rect -5036 -3000 -4996 -1680
rect -6396 -3040 -4996 -3000
rect -3898 -1680 -2498 -1640
rect -3898 -3000 -3858 -1680
rect -2538 -3000 -2498 -1680
rect -3898 -3040 -2498 -3000
rect -1400 -1680 0 -1640
rect -1400 -3000 -1360 -1680
rect -40 -3000 0 -1680
rect -1400 -3040 0 -3000
rect 1098 -1680 2498 -1640
rect 1098 -3000 1138 -1680
rect 2458 -3000 2498 -1680
rect 1098 -3040 2498 -3000
rect 3596 -1680 4996 -1640
rect 3596 -3000 3636 -1680
rect 4956 -3000 4996 -1680
rect 3596 -3040 4996 -3000
rect 6094 -1680 7494 -1640
rect 6094 -3000 6134 -1680
rect 7454 -3000 7494 -1680
rect 6094 -3040 7494 -3000
rect 8592 -1680 9992 -1640
rect 8592 -3000 8632 -1680
rect 9952 -3000 9992 -1680
rect 8592 -3040 9992 -3000
rect 11090 -1680 12490 -1640
rect 11090 -3000 11130 -1680
rect 12450 -3000 12490 -1680
rect 11090 -3040 12490 -3000
rect -8894 -3480 -7494 -3440
rect -8894 -4800 -8854 -3480
rect -7534 -4800 -7494 -3480
rect -8894 -4840 -7494 -4800
rect -6396 -3480 -4996 -3440
rect -6396 -4800 -6356 -3480
rect -5036 -4800 -4996 -3480
rect -6396 -4840 -4996 -4800
rect -3898 -3480 -2498 -3440
rect -3898 -4800 -3858 -3480
rect -2538 -4800 -2498 -3480
rect -3898 -4840 -2498 -4800
rect -1400 -3480 0 -3440
rect -1400 -4800 -1360 -3480
rect -40 -4800 0 -3480
rect -1400 -4840 0 -4800
rect 1098 -3480 2498 -3440
rect 1098 -4800 1138 -3480
rect 2458 -4800 2498 -3480
rect 1098 -4840 2498 -4800
rect 3596 -3480 4996 -3440
rect 3596 -4800 3636 -3480
rect 4956 -4800 4996 -3480
rect 3596 -4840 4996 -4800
rect 6094 -3480 7494 -3440
rect 6094 -4800 6134 -3480
rect 7454 -4800 7494 -3480
rect 6094 -4840 7494 -4800
rect 8592 -3480 9992 -3440
rect 8592 -4800 8632 -3480
rect 9952 -4800 9992 -3480
rect 8592 -4840 9992 -4800
rect 11090 -3480 12490 -3440
rect 11090 -4800 11130 -3480
rect 12450 -4800 12490 -3480
rect 11090 -4840 12490 -4800
rect -8894 -5280 -7494 -5240
rect -8894 -6600 -8854 -5280
rect -7534 -6600 -7494 -5280
rect -8894 -6640 -7494 -6600
rect -6396 -5280 -4996 -5240
rect -6396 -6600 -6356 -5280
rect -5036 -6600 -4996 -5280
rect -6396 -6640 -4996 -6600
rect -3898 -5280 -2498 -5240
rect -3898 -6600 -3858 -5280
rect -2538 -6600 -2498 -5280
rect -3898 -6640 -2498 -6600
rect -1400 -5280 0 -5240
rect -1400 -6600 -1360 -5280
rect -40 -6600 0 -5280
rect -1400 -6640 0 -6600
rect 1098 -5280 2498 -5240
rect 1098 -6600 1138 -5280
rect 2458 -6600 2498 -5280
rect 1098 -6640 2498 -6600
rect 3596 -5280 4996 -5240
rect 3596 -6600 3636 -5280
rect 4956 -6600 4996 -5280
rect 3596 -6640 4996 -6600
rect 6094 -5280 7494 -5240
rect 6094 -6600 6134 -5280
rect 7454 -6600 7494 -5280
rect 6094 -6640 7494 -6600
rect 8592 -5280 9992 -5240
rect 8592 -6600 8632 -5280
rect 9952 -6600 9992 -5280
rect 8592 -6640 9992 -6600
rect 11090 -5280 12490 -5240
rect 11090 -6600 11130 -5280
rect 12450 -6600 12490 -5280
rect 11090 -6640 12490 -6600
rect -8894 -7080 -7494 -7040
rect -8894 -8400 -8854 -7080
rect -7534 -8400 -7494 -7080
rect -8894 -8440 -7494 -8400
rect -6396 -7080 -4996 -7040
rect -6396 -8400 -6356 -7080
rect -5036 -8400 -4996 -7080
rect -6396 -8440 -4996 -8400
rect -3898 -7080 -2498 -7040
rect -3898 -8400 -3858 -7080
rect -2538 -8400 -2498 -7080
rect -3898 -8440 -2498 -8400
rect -1400 -7080 0 -7040
rect -1400 -8400 -1360 -7080
rect -40 -8400 0 -7080
rect -1400 -8440 0 -8400
rect 1098 -7080 2498 -7040
rect 1098 -8400 1138 -7080
rect 2458 -8400 2498 -7080
rect 1098 -8440 2498 -8400
rect 3596 -7080 4996 -7040
rect 3596 -8400 3636 -7080
rect 4956 -8400 4996 -7080
rect 3596 -8440 4996 -8400
rect 6094 -7080 7494 -7040
rect 6094 -8400 6134 -7080
rect 7454 -8400 7494 -7080
rect 6094 -8440 7494 -8400
rect 8592 -7080 9992 -7040
rect 8592 -8400 8632 -7080
rect 9952 -8400 9992 -7080
rect 8592 -8440 9992 -8400
rect 11090 -7080 12490 -7040
rect 11090 -8400 11130 -7080
rect 12450 -8400 12490 -7080
rect 11090 -8440 12490 -8400
<< mimcapcontact >>
rect -8854 7800 -7534 9120
rect -6356 7800 -5036 9120
rect -3858 7800 -2538 9120
rect -1360 7800 -40 9120
rect 1138 7800 2458 9120
rect 3636 7800 4956 9120
rect 6134 7800 7454 9120
rect 8632 7800 9952 9120
rect 11130 7800 12450 9120
rect -8854 6000 -7534 7320
rect -6356 6000 -5036 7320
rect -3858 6000 -2538 7320
rect -1360 6000 -40 7320
rect 1138 6000 2458 7320
rect 3636 6000 4956 7320
rect 6134 6000 7454 7320
rect 8632 6000 9952 7320
rect 11130 6000 12450 7320
rect -8854 4200 -7534 5520
rect -6356 4200 -5036 5520
rect -3858 4200 -2538 5520
rect -1360 4200 -40 5520
rect 1138 4200 2458 5520
rect 3636 4200 4956 5520
rect 6134 4200 7454 5520
rect 8632 4200 9952 5520
rect 11130 4200 12450 5520
rect -8854 2400 -7534 3720
rect -6356 2400 -5036 3720
rect -3858 2400 -2538 3720
rect -1360 2400 -40 3720
rect 1138 2400 2458 3720
rect 3636 2400 4956 3720
rect 6134 2400 7454 3720
rect 8632 2400 9952 3720
rect 11130 2400 12450 3720
rect -8854 600 -7534 1920
rect -6356 600 -5036 1920
rect -3858 600 -2538 1920
rect -1360 600 -40 1920
rect 1138 600 2458 1920
rect 3636 600 4956 1920
rect 6134 600 7454 1920
rect 8632 600 9952 1920
rect 11130 600 12450 1920
rect -8854 -1200 -7534 120
rect -6356 -1200 -5036 120
rect -3858 -1200 -2538 120
rect -1360 -1200 -40 120
rect 1138 -1200 2458 120
rect 3636 -1200 4956 120
rect 6134 -1200 7454 120
rect 8632 -1200 9952 120
rect 11130 -1200 12450 120
rect -8854 -3000 -7534 -1680
rect -6356 -3000 -5036 -1680
rect -3858 -3000 -2538 -1680
rect -1360 -3000 -40 -1680
rect 1138 -3000 2458 -1680
rect 3636 -3000 4956 -1680
rect 6134 -3000 7454 -1680
rect 8632 -3000 9952 -1680
rect 11130 -3000 12450 -1680
rect -8854 -4800 -7534 -3480
rect -6356 -4800 -5036 -3480
rect -3858 -4800 -2538 -3480
rect -1360 -4800 -40 -3480
rect 1138 -4800 2458 -3480
rect 3636 -4800 4956 -3480
rect 6134 -4800 7454 -3480
rect 8632 -4800 9952 -3480
rect 11130 -4800 12450 -3480
rect -8854 -6600 -7534 -5280
rect -6356 -6600 -5036 -5280
rect -3858 -6600 -2538 -5280
rect -1360 -6600 -40 -5280
rect 1138 -6600 2458 -5280
rect 3636 -6600 4956 -5280
rect 6134 -6600 7454 -5280
rect 8632 -6600 9952 -5280
rect 11130 -6600 12450 -5280
rect -8854 -8400 -7534 -7080
rect -6356 -8400 -5036 -7080
rect -3858 -8400 -2538 -7080
rect -1360 -8400 -40 -7080
rect 1138 -8400 2458 -7080
rect 3636 -8400 4956 -7080
rect 6134 -8400 7454 -7080
rect 8632 -8400 9952 -7080
rect 11130 -8400 12450 -7080
<< metal4 >>
rect -7262 9172 -7166 9188
rect -8855 9120 -7533 9121
rect -8855 7800 -8854 9120
rect -7534 7800 -7533 9120
rect -8855 7799 -7533 7800
rect -7262 7748 -7246 9172
rect -7182 7748 -7166 9172
rect -4764 9172 -4668 9188
rect -6357 9120 -5035 9121
rect -6357 7800 -6356 9120
rect -5036 7800 -5035 9120
rect -6357 7799 -5035 7800
rect -7262 7732 -7166 7748
rect -4764 7748 -4748 9172
rect -4684 7748 -4668 9172
rect -2266 9172 -2170 9188
rect -3859 9120 -2537 9121
rect -3859 7800 -3858 9120
rect -2538 7800 -2537 9120
rect -3859 7799 -2537 7800
rect -4764 7732 -4668 7748
rect -2266 7748 -2250 9172
rect -2186 7748 -2170 9172
rect 232 9172 328 9188
rect -1361 9120 -39 9121
rect -1361 7800 -1360 9120
rect -40 7800 -39 9120
rect -1361 7799 -39 7800
rect -2266 7732 -2170 7748
rect 232 7748 248 9172
rect 312 7748 328 9172
rect 2730 9172 2826 9188
rect 1137 9120 2459 9121
rect 1137 7800 1138 9120
rect 2458 7800 2459 9120
rect 1137 7799 2459 7800
rect 232 7732 328 7748
rect 2730 7748 2746 9172
rect 2810 7748 2826 9172
rect 5228 9172 5324 9188
rect 3635 9120 4957 9121
rect 3635 7800 3636 9120
rect 4956 7800 4957 9120
rect 3635 7799 4957 7800
rect 2730 7732 2826 7748
rect 5228 7748 5244 9172
rect 5308 7748 5324 9172
rect 7726 9172 7822 9188
rect 6133 9120 7455 9121
rect 6133 7800 6134 9120
rect 7454 7800 7455 9120
rect 6133 7799 7455 7800
rect 5228 7732 5324 7748
rect 7726 7748 7742 9172
rect 7806 7748 7822 9172
rect 10224 9172 10320 9188
rect 8631 9120 9953 9121
rect 8631 7800 8632 9120
rect 9952 7800 9953 9120
rect 8631 7799 9953 7800
rect 7726 7732 7822 7748
rect 10224 7748 10240 9172
rect 10304 7748 10320 9172
rect 12722 9172 12818 9188
rect 11129 9120 12451 9121
rect 11129 7800 11130 9120
rect 12450 7800 12451 9120
rect 11129 7799 12451 7800
rect 10224 7732 10320 7748
rect 12722 7748 12738 9172
rect 12802 7748 12818 9172
rect 12722 7732 12818 7748
rect -7262 7372 -7166 7388
rect -8855 7320 -7533 7321
rect -8855 6000 -8854 7320
rect -7534 6000 -7533 7320
rect -8855 5999 -7533 6000
rect -7262 5948 -7246 7372
rect -7182 5948 -7166 7372
rect -4764 7372 -4668 7388
rect -6357 7320 -5035 7321
rect -6357 6000 -6356 7320
rect -5036 6000 -5035 7320
rect -6357 5999 -5035 6000
rect -7262 5932 -7166 5948
rect -4764 5948 -4748 7372
rect -4684 5948 -4668 7372
rect -2266 7372 -2170 7388
rect -3859 7320 -2537 7321
rect -3859 6000 -3858 7320
rect -2538 6000 -2537 7320
rect -3859 5999 -2537 6000
rect -4764 5932 -4668 5948
rect -2266 5948 -2250 7372
rect -2186 5948 -2170 7372
rect 232 7372 328 7388
rect -1361 7320 -39 7321
rect -1361 6000 -1360 7320
rect -40 6000 -39 7320
rect -1361 5999 -39 6000
rect -2266 5932 -2170 5948
rect 232 5948 248 7372
rect 312 5948 328 7372
rect 2730 7372 2826 7388
rect 1137 7320 2459 7321
rect 1137 6000 1138 7320
rect 2458 6000 2459 7320
rect 1137 5999 2459 6000
rect 232 5932 328 5948
rect 2730 5948 2746 7372
rect 2810 5948 2826 7372
rect 5228 7372 5324 7388
rect 3635 7320 4957 7321
rect 3635 6000 3636 7320
rect 4956 6000 4957 7320
rect 3635 5999 4957 6000
rect 2730 5932 2826 5948
rect 5228 5948 5244 7372
rect 5308 5948 5324 7372
rect 7726 7372 7822 7388
rect 6133 7320 7455 7321
rect 6133 6000 6134 7320
rect 7454 6000 7455 7320
rect 6133 5999 7455 6000
rect 5228 5932 5324 5948
rect 7726 5948 7742 7372
rect 7806 5948 7822 7372
rect 10224 7372 10320 7388
rect 8631 7320 9953 7321
rect 8631 6000 8632 7320
rect 9952 6000 9953 7320
rect 8631 5999 9953 6000
rect 7726 5932 7822 5948
rect 10224 5948 10240 7372
rect 10304 5948 10320 7372
rect 12722 7372 12818 7388
rect 11129 7320 12451 7321
rect 11129 6000 11130 7320
rect 12450 6000 12451 7320
rect 11129 5999 12451 6000
rect 10224 5932 10320 5948
rect 12722 5948 12738 7372
rect 12802 5948 12818 7372
rect 12722 5932 12818 5948
rect -7262 5572 -7166 5588
rect -8855 5520 -7533 5521
rect -8855 4200 -8854 5520
rect -7534 4200 -7533 5520
rect -8855 4199 -7533 4200
rect -7262 4148 -7246 5572
rect -7182 4148 -7166 5572
rect -4764 5572 -4668 5588
rect -6357 5520 -5035 5521
rect -6357 4200 -6356 5520
rect -5036 4200 -5035 5520
rect -6357 4199 -5035 4200
rect -7262 4132 -7166 4148
rect -4764 4148 -4748 5572
rect -4684 4148 -4668 5572
rect -2266 5572 -2170 5588
rect -3859 5520 -2537 5521
rect -3859 4200 -3858 5520
rect -2538 4200 -2537 5520
rect -3859 4199 -2537 4200
rect -4764 4132 -4668 4148
rect -2266 4148 -2250 5572
rect -2186 4148 -2170 5572
rect 232 5572 328 5588
rect -1361 5520 -39 5521
rect -1361 4200 -1360 5520
rect -40 4200 -39 5520
rect -1361 4199 -39 4200
rect -2266 4132 -2170 4148
rect 232 4148 248 5572
rect 312 4148 328 5572
rect 2730 5572 2826 5588
rect 1137 5520 2459 5521
rect 1137 4200 1138 5520
rect 2458 4200 2459 5520
rect 1137 4199 2459 4200
rect 232 4132 328 4148
rect 2730 4148 2746 5572
rect 2810 4148 2826 5572
rect 5228 5572 5324 5588
rect 3635 5520 4957 5521
rect 3635 4200 3636 5520
rect 4956 4200 4957 5520
rect 3635 4199 4957 4200
rect 2730 4132 2826 4148
rect 5228 4148 5244 5572
rect 5308 4148 5324 5572
rect 7726 5572 7822 5588
rect 6133 5520 7455 5521
rect 6133 4200 6134 5520
rect 7454 4200 7455 5520
rect 6133 4199 7455 4200
rect 5228 4132 5324 4148
rect 7726 4148 7742 5572
rect 7806 4148 7822 5572
rect 10224 5572 10320 5588
rect 8631 5520 9953 5521
rect 8631 4200 8632 5520
rect 9952 4200 9953 5520
rect 8631 4199 9953 4200
rect 7726 4132 7822 4148
rect 10224 4148 10240 5572
rect 10304 4148 10320 5572
rect 12722 5572 12818 5588
rect 11129 5520 12451 5521
rect 11129 4200 11130 5520
rect 12450 4200 12451 5520
rect 11129 4199 12451 4200
rect 10224 4132 10320 4148
rect 12722 4148 12738 5572
rect 12802 4148 12818 5572
rect 12722 4132 12818 4148
rect -7262 3772 -7166 3788
rect -8855 3720 -7533 3721
rect -8855 2400 -8854 3720
rect -7534 2400 -7533 3720
rect -8855 2399 -7533 2400
rect -7262 2348 -7246 3772
rect -7182 2348 -7166 3772
rect -4764 3772 -4668 3788
rect -6357 3720 -5035 3721
rect -6357 2400 -6356 3720
rect -5036 2400 -5035 3720
rect -6357 2399 -5035 2400
rect -7262 2332 -7166 2348
rect -4764 2348 -4748 3772
rect -4684 2348 -4668 3772
rect -2266 3772 -2170 3788
rect -3859 3720 -2537 3721
rect -3859 2400 -3858 3720
rect -2538 2400 -2537 3720
rect -3859 2399 -2537 2400
rect -4764 2332 -4668 2348
rect -2266 2348 -2250 3772
rect -2186 2348 -2170 3772
rect 232 3772 328 3788
rect -1361 3720 -39 3721
rect -1361 2400 -1360 3720
rect -40 2400 -39 3720
rect -1361 2399 -39 2400
rect -2266 2332 -2170 2348
rect 232 2348 248 3772
rect 312 2348 328 3772
rect 2730 3772 2826 3788
rect 1137 3720 2459 3721
rect 1137 2400 1138 3720
rect 2458 2400 2459 3720
rect 1137 2399 2459 2400
rect 232 2332 328 2348
rect 2730 2348 2746 3772
rect 2810 2348 2826 3772
rect 5228 3772 5324 3788
rect 3635 3720 4957 3721
rect 3635 2400 3636 3720
rect 4956 2400 4957 3720
rect 3635 2399 4957 2400
rect 2730 2332 2826 2348
rect 5228 2348 5244 3772
rect 5308 2348 5324 3772
rect 7726 3772 7822 3788
rect 6133 3720 7455 3721
rect 6133 2400 6134 3720
rect 7454 2400 7455 3720
rect 6133 2399 7455 2400
rect 5228 2332 5324 2348
rect 7726 2348 7742 3772
rect 7806 2348 7822 3772
rect 10224 3772 10320 3788
rect 8631 3720 9953 3721
rect 8631 2400 8632 3720
rect 9952 2400 9953 3720
rect 8631 2399 9953 2400
rect 7726 2332 7822 2348
rect 10224 2348 10240 3772
rect 10304 2348 10320 3772
rect 12722 3772 12818 3788
rect 11129 3720 12451 3721
rect 11129 2400 11130 3720
rect 12450 2400 12451 3720
rect 11129 2399 12451 2400
rect 10224 2332 10320 2348
rect 12722 2348 12738 3772
rect 12802 2348 12818 3772
rect 12722 2332 12818 2348
rect -7262 1972 -7166 1988
rect -8855 1920 -7533 1921
rect -8855 600 -8854 1920
rect -7534 600 -7533 1920
rect -8855 599 -7533 600
rect -7262 548 -7246 1972
rect -7182 548 -7166 1972
rect -4764 1972 -4668 1988
rect -6357 1920 -5035 1921
rect -6357 600 -6356 1920
rect -5036 600 -5035 1920
rect -6357 599 -5035 600
rect -7262 532 -7166 548
rect -4764 548 -4748 1972
rect -4684 548 -4668 1972
rect -2266 1972 -2170 1988
rect -3859 1920 -2537 1921
rect -3859 600 -3858 1920
rect -2538 600 -2537 1920
rect -3859 599 -2537 600
rect -4764 532 -4668 548
rect -2266 548 -2250 1972
rect -2186 548 -2170 1972
rect 232 1972 328 1988
rect -1361 1920 -39 1921
rect -1361 600 -1360 1920
rect -40 600 -39 1920
rect -1361 599 -39 600
rect -2266 532 -2170 548
rect 232 548 248 1972
rect 312 548 328 1972
rect 2730 1972 2826 1988
rect 1137 1920 2459 1921
rect 1137 600 1138 1920
rect 2458 600 2459 1920
rect 1137 599 2459 600
rect 232 532 328 548
rect 2730 548 2746 1972
rect 2810 548 2826 1972
rect 5228 1972 5324 1988
rect 3635 1920 4957 1921
rect 3635 600 3636 1920
rect 4956 600 4957 1920
rect 3635 599 4957 600
rect 2730 532 2826 548
rect 5228 548 5244 1972
rect 5308 548 5324 1972
rect 7726 1972 7822 1988
rect 6133 1920 7455 1921
rect 6133 600 6134 1920
rect 7454 600 7455 1920
rect 6133 599 7455 600
rect 5228 532 5324 548
rect 7726 548 7742 1972
rect 7806 548 7822 1972
rect 10224 1972 10320 1988
rect 8631 1920 9953 1921
rect 8631 600 8632 1920
rect 9952 600 9953 1920
rect 8631 599 9953 600
rect 7726 532 7822 548
rect 10224 548 10240 1972
rect 10304 548 10320 1972
rect 12722 1972 12818 1988
rect 11129 1920 12451 1921
rect 11129 600 11130 1920
rect 12450 600 12451 1920
rect 11129 599 12451 600
rect 10224 532 10320 548
rect 12722 548 12738 1972
rect 12802 548 12818 1972
rect 12722 532 12818 548
rect -7262 172 -7166 188
rect -8855 120 -7533 121
rect -8855 -1200 -8854 120
rect -7534 -1200 -7533 120
rect -8855 -1201 -7533 -1200
rect -7262 -1252 -7246 172
rect -7182 -1252 -7166 172
rect -4764 172 -4668 188
rect -6357 120 -5035 121
rect -6357 -1200 -6356 120
rect -5036 -1200 -5035 120
rect -6357 -1201 -5035 -1200
rect -7262 -1268 -7166 -1252
rect -4764 -1252 -4748 172
rect -4684 -1252 -4668 172
rect -2266 172 -2170 188
rect -3859 120 -2537 121
rect -3859 -1200 -3858 120
rect -2538 -1200 -2537 120
rect -3859 -1201 -2537 -1200
rect -4764 -1268 -4668 -1252
rect -2266 -1252 -2250 172
rect -2186 -1252 -2170 172
rect 232 172 328 188
rect -1361 120 -39 121
rect -1361 -1200 -1360 120
rect -40 -1200 -39 120
rect -1361 -1201 -39 -1200
rect -2266 -1268 -2170 -1252
rect 232 -1252 248 172
rect 312 -1252 328 172
rect 2730 172 2826 188
rect 1137 120 2459 121
rect 1137 -1200 1138 120
rect 2458 -1200 2459 120
rect 1137 -1201 2459 -1200
rect 232 -1268 328 -1252
rect 2730 -1252 2746 172
rect 2810 -1252 2826 172
rect 5228 172 5324 188
rect 3635 120 4957 121
rect 3635 -1200 3636 120
rect 4956 -1200 4957 120
rect 3635 -1201 4957 -1200
rect 2730 -1268 2826 -1252
rect 5228 -1252 5244 172
rect 5308 -1252 5324 172
rect 7726 172 7822 188
rect 6133 120 7455 121
rect 6133 -1200 6134 120
rect 7454 -1200 7455 120
rect 6133 -1201 7455 -1200
rect 5228 -1268 5324 -1252
rect 7726 -1252 7742 172
rect 7806 -1252 7822 172
rect 10224 172 10320 188
rect 8631 120 9953 121
rect 8631 -1200 8632 120
rect 9952 -1200 9953 120
rect 8631 -1201 9953 -1200
rect 7726 -1268 7822 -1252
rect 10224 -1252 10240 172
rect 10304 -1252 10320 172
rect 12722 172 12818 188
rect 11129 120 12451 121
rect 11129 -1200 11130 120
rect 12450 -1200 12451 120
rect 11129 -1201 12451 -1200
rect 10224 -1268 10320 -1252
rect 12722 -1252 12738 172
rect 12802 -1252 12818 172
rect 12722 -1268 12818 -1252
rect -7262 -1628 -7166 -1612
rect -8855 -1680 -7533 -1679
rect -8855 -3000 -8854 -1680
rect -7534 -3000 -7533 -1680
rect -8855 -3001 -7533 -3000
rect -7262 -3052 -7246 -1628
rect -7182 -3052 -7166 -1628
rect -4764 -1628 -4668 -1612
rect -6357 -1680 -5035 -1679
rect -6357 -3000 -6356 -1680
rect -5036 -3000 -5035 -1680
rect -6357 -3001 -5035 -3000
rect -7262 -3068 -7166 -3052
rect -4764 -3052 -4748 -1628
rect -4684 -3052 -4668 -1628
rect -2266 -1628 -2170 -1612
rect -3859 -1680 -2537 -1679
rect -3859 -3000 -3858 -1680
rect -2538 -3000 -2537 -1680
rect -3859 -3001 -2537 -3000
rect -4764 -3068 -4668 -3052
rect -2266 -3052 -2250 -1628
rect -2186 -3052 -2170 -1628
rect 232 -1628 328 -1612
rect -1361 -1680 -39 -1679
rect -1361 -3000 -1360 -1680
rect -40 -3000 -39 -1680
rect -1361 -3001 -39 -3000
rect -2266 -3068 -2170 -3052
rect 232 -3052 248 -1628
rect 312 -3052 328 -1628
rect 2730 -1628 2826 -1612
rect 1137 -1680 2459 -1679
rect 1137 -3000 1138 -1680
rect 2458 -3000 2459 -1680
rect 1137 -3001 2459 -3000
rect 232 -3068 328 -3052
rect 2730 -3052 2746 -1628
rect 2810 -3052 2826 -1628
rect 5228 -1628 5324 -1612
rect 3635 -1680 4957 -1679
rect 3635 -3000 3636 -1680
rect 4956 -3000 4957 -1680
rect 3635 -3001 4957 -3000
rect 2730 -3068 2826 -3052
rect 5228 -3052 5244 -1628
rect 5308 -3052 5324 -1628
rect 7726 -1628 7822 -1612
rect 6133 -1680 7455 -1679
rect 6133 -3000 6134 -1680
rect 7454 -3000 7455 -1680
rect 6133 -3001 7455 -3000
rect 5228 -3068 5324 -3052
rect 7726 -3052 7742 -1628
rect 7806 -3052 7822 -1628
rect 10224 -1628 10320 -1612
rect 8631 -1680 9953 -1679
rect 8631 -3000 8632 -1680
rect 9952 -3000 9953 -1680
rect 8631 -3001 9953 -3000
rect 7726 -3068 7822 -3052
rect 10224 -3052 10240 -1628
rect 10304 -3052 10320 -1628
rect 12722 -1628 12818 -1612
rect 11129 -1680 12451 -1679
rect 11129 -3000 11130 -1680
rect 12450 -3000 12451 -1680
rect 11129 -3001 12451 -3000
rect 10224 -3068 10320 -3052
rect 12722 -3052 12738 -1628
rect 12802 -3052 12818 -1628
rect 12722 -3068 12818 -3052
rect -7262 -3428 -7166 -3412
rect -8855 -3480 -7533 -3479
rect -8855 -4800 -8854 -3480
rect -7534 -4800 -7533 -3480
rect -8855 -4801 -7533 -4800
rect -7262 -4852 -7246 -3428
rect -7182 -4852 -7166 -3428
rect -4764 -3428 -4668 -3412
rect -6357 -3480 -5035 -3479
rect -6357 -4800 -6356 -3480
rect -5036 -4800 -5035 -3480
rect -6357 -4801 -5035 -4800
rect -7262 -4868 -7166 -4852
rect -4764 -4852 -4748 -3428
rect -4684 -4852 -4668 -3428
rect -2266 -3428 -2170 -3412
rect -3859 -3480 -2537 -3479
rect -3859 -4800 -3858 -3480
rect -2538 -4800 -2537 -3480
rect -3859 -4801 -2537 -4800
rect -4764 -4868 -4668 -4852
rect -2266 -4852 -2250 -3428
rect -2186 -4852 -2170 -3428
rect 232 -3428 328 -3412
rect -1361 -3480 -39 -3479
rect -1361 -4800 -1360 -3480
rect -40 -4800 -39 -3480
rect -1361 -4801 -39 -4800
rect -2266 -4868 -2170 -4852
rect 232 -4852 248 -3428
rect 312 -4852 328 -3428
rect 2730 -3428 2826 -3412
rect 1137 -3480 2459 -3479
rect 1137 -4800 1138 -3480
rect 2458 -4800 2459 -3480
rect 1137 -4801 2459 -4800
rect 232 -4868 328 -4852
rect 2730 -4852 2746 -3428
rect 2810 -4852 2826 -3428
rect 5228 -3428 5324 -3412
rect 3635 -3480 4957 -3479
rect 3635 -4800 3636 -3480
rect 4956 -4800 4957 -3480
rect 3635 -4801 4957 -4800
rect 2730 -4868 2826 -4852
rect 5228 -4852 5244 -3428
rect 5308 -4852 5324 -3428
rect 7726 -3428 7822 -3412
rect 6133 -3480 7455 -3479
rect 6133 -4800 6134 -3480
rect 7454 -4800 7455 -3480
rect 6133 -4801 7455 -4800
rect 5228 -4868 5324 -4852
rect 7726 -4852 7742 -3428
rect 7806 -4852 7822 -3428
rect 10224 -3428 10320 -3412
rect 8631 -3480 9953 -3479
rect 8631 -4800 8632 -3480
rect 9952 -4800 9953 -3480
rect 8631 -4801 9953 -4800
rect 7726 -4868 7822 -4852
rect 10224 -4852 10240 -3428
rect 10304 -4852 10320 -3428
rect 12722 -3428 12818 -3412
rect 11129 -3480 12451 -3479
rect 11129 -4800 11130 -3480
rect 12450 -4800 12451 -3480
rect 11129 -4801 12451 -4800
rect 10224 -4868 10320 -4852
rect 12722 -4852 12738 -3428
rect 12802 -4852 12818 -3428
rect 12722 -4868 12818 -4852
rect -7262 -5228 -7166 -5212
rect -8855 -5280 -7533 -5279
rect -8855 -6600 -8854 -5280
rect -7534 -6600 -7533 -5280
rect -8855 -6601 -7533 -6600
rect -7262 -6652 -7246 -5228
rect -7182 -6652 -7166 -5228
rect -4764 -5228 -4668 -5212
rect -6357 -5280 -5035 -5279
rect -6357 -6600 -6356 -5280
rect -5036 -6600 -5035 -5280
rect -6357 -6601 -5035 -6600
rect -7262 -6668 -7166 -6652
rect -4764 -6652 -4748 -5228
rect -4684 -6652 -4668 -5228
rect -2266 -5228 -2170 -5212
rect -3859 -5280 -2537 -5279
rect -3859 -6600 -3858 -5280
rect -2538 -6600 -2537 -5280
rect -3859 -6601 -2537 -6600
rect -4764 -6668 -4668 -6652
rect -2266 -6652 -2250 -5228
rect -2186 -6652 -2170 -5228
rect 232 -5228 328 -5212
rect -1361 -5280 -39 -5279
rect -1361 -6600 -1360 -5280
rect -40 -6600 -39 -5280
rect -1361 -6601 -39 -6600
rect -2266 -6668 -2170 -6652
rect 232 -6652 248 -5228
rect 312 -6652 328 -5228
rect 2730 -5228 2826 -5212
rect 1137 -5280 2459 -5279
rect 1137 -6600 1138 -5280
rect 2458 -6600 2459 -5280
rect 1137 -6601 2459 -6600
rect 232 -6668 328 -6652
rect 2730 -6652 2746 -5228
rect 2810 -6652 2826 -5228
rect 5228 -5228 5324 -5212
rect 3635 -5280 4957 -5279
rect 3635 -6600 3636 -5280
rect 4956 -6600 4957 -5280
rect 3635 -6601 4957 -6600
rect 2730 -6668 2826 -6652
rect 5228 -6652 5244 -5228
rect 5308 -6652 5324 -5228
rect 7726 -5228 7822 -5212
rect 6133 -5280 7455 -5279
rect 6133 -6600 6134 -5280
rect 7454 -6600 7455 -5280
rect 6133 -6601 7455 -6600
rect 5228 -6668 5324 -6652
rect 7726 -6652 7742 -5228
rect 7806 -6652 7822 -5228
rect 10224 -5228 10320 -5212
rect 8631 -5280 9953 -5279
rect 8631 -6600 8632 -5280
rect 9952 -6600 9953 -5280
rect 8631 -6601 9953 -6600
rect 7726 -6668 7822 -6652
rect 10224 -6652 10240 -5228
rect 10304 -6652 10320 -5228
rect 12722 -5228 12818 -5212
rect 11129 -5280 12451 -5279
rect 11129 -6600 11130 -5280
rect 12450 -6600 12451 -5280
rect 11129 -6601 12451 -6600
rect 10224 -6668 10320 -6652
rect 12722 -6652 12738 -5228
rect 12802 -6652 12818 -5228
rect 12722 -6668 12818 -6652
rect -7262 -7028 -7166 -7012
rect -8855 -7080 -7533 -7079
rect -8855 -8400 -8854 -7080
rect -7534 -8400 -7533 -7080
rect -8855 -8401 -7533 -8400
rect -7262 -8452 -7246 -7028
rect -7182 -8452 -7166 -7028
rect -4764 -7028 -4668 -7012
rect -6357 -7080 -5035 -7079
rect -6357 -8400 -6356 -7080
rect -5036 -8400 -5035 -7080
rect -6357 -8401 -5035 -8400
rect -7262 -8468 -7166 -8452
rect -4764 -8452 -4748 -7028
rect -4684 -8452 -4668 -7028
rect -2266 -7028 -2170 -7012
rect -3859 -7080 -2537 -7079
rect -3859 -8400 -3858 -7080
rect -2538 -8400 -2537 -7080
rect -3859 -8401 -2537 -8400
rect -4764 -8468 -4668 -8452
rect -2266 -8452 -2250 -7028
rect -2186 -8452 -2170 -7028
rect 232 -7028 328 -7012
rect -1361 -7080 -39 -7079
rect -1361 -8400 -1360 -7080
rect -40 -8400 -39 -7080
rect -1361 -8401 -39 -8400
rect -2266 -8468 -2170 -8452
rect 232 -8452 248 -7028
rect 312 -8452 328 -7028
rect 2730 -7028 2826 -7012
rect 1137 -7080 2459 -7079
rect 1137 -8400 1138 -7080
rect 2458 -8400 2459 -7080
rect 1137 -8401 2459 -8400
rect 232 -8468 328 -8452
rect 2730 -8452 2746 -7028
rect 2810 -8452 2826 -7028
rect 5228 -7028 5324 -7012
rect 3635 -7080 4957 -7079
rect 3635 -8400 3636 -7080
rect 4956 -8400 4957 -7080
rect 3635 -8401 4957 -8400
rect 2730 -8468 2826 -8452
rect 5228 -8452 5244 -7028
rect 5308 -8452 5324 -7028
rect 7726 -7028 7822 -7012
rect 6133 -7080 7455 -7079
rect 6133 -8400 6134 -7080
rect 7454 -8400 7455 -7080
rect 6133 -8401 7455 -8400
rect 5228 -8468 5324 -8452
rect 7726 -8452 7742 -7028
rect 7806 -8452 7822 -7028
rect 10224 -7028 10320 -7012
rect 8631 -7080 9953 -7079
rect 8631 -8400 8632 -7080
rect 9952 -8400 9953 -7080
rect 8631 -8401 9953 -8400
rect 7726 -8468 7822 -8452
rect 10224 -8452 10240 -7028
rect 10304 -8452 10320 -7028
rect 12722 -7028 12818 -7012
rect 11129 -7080 12451 -7079
rect 11129 -8400 11130 -7080
rect 12450 -8400 12451 -7080
rect 11129 -8401 12451 -8400
rect 10224 -8468 10320 -8452
rect 12722 -8452 12738 -7028
rect 12802 -8452 12818 -7028
rect 12722 -8468 12818 -8452
<< properties >>
string FIXED_BBOX 7162 7000 8642 8480
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7.0 l 7.0 val 103.32 carea 2.00 cperi 0.19 nx 9 ny 10 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
