** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/sky130_ef_ip__cdac3v_12bit.sch
.subckt sky130_ef_ip__cdac3v_12bit SELD0 SELD1 SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8 SELD9 VDD DVDD DVSS VSS VH VL OUT RST
+ OUTNC SELD10 SELD11
*.PININFO SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VDD:B DVDD:B DVSS:B VH:B VL:B VSS:B
*+ RST:I OUT:O OUTNC:O SELD10:I SELD11:I
x4 D8 D0 D4 OUTNC D9 D5 D1 OUT D2 D6 VSS D7 D3 D10 D11 EF_BANK_CAP_12
x3 D0 SELD0 D1 SELD1 SELD2 D2 SELD3 SELD4 D3 SELD5 D4 SELD6 SELD7 D5 SELD8 D6 SELD9 D7 D8 D9 VDD DVDD DVSS VH VL VSS D10 D11
+ SELD10 SELD11 EF_AMUX0201_ARRAY1
x1 OUTNC OUT VDD DVDD VSS RST DVSS EF_SW_RST
.ends

* expanding   symbol:  EF_BANK_CAP_12.sym # of pins=15
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_BANK_CAP_12.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_BANK_CAP_12.sch
.subckt EF_BANK_CAP_12 D8 D0 D4 VP1 D9 D5 D1 VP2 D2 D6 VSS D7 D3 D10 D11
*.PININFO D0:B D1:B D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B VSS:B VP1:B VP2:B D10:B D11:B
x4 VP1 VSS D0 D1 D2 D3 D4 D5 EF_LSB_CAP
x1 D8 D10 D9 VP2 D6 VSS D7 D11 EF_MSB_CAP
x2 VP1 VP2 VSS EF_SC_CAP
.ends


* expanding   symbol:  EF_AMUX0201_ARRAY1.sym # of pins=30
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX0201_ARRAY1.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX0201_ARRAY1.sch
.subckt EF_AMUX0201_ARRAY1 D0 SELD0 D1 SELD1 SELD2 D2 SELD3 SELD4 D3 SELD5 D4 SELD6 SELD7 D5 SELD8 D6 SELD9 D7 D8 D9 VDD DVDD DVSS
+ VH VL VSS D10 D11 SELD10 SELD11
*.PININFO VDD:B DVDD:B DVSS:B VH:B VL:B SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VSS:B D0:B
*+ D1:B D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B SELD10:I SELD11:I D10:B D11:B
x2 VDD DVDD D0 VSS VH VL SELD0 DVSS EF_AMUX21x
x1 VDD DVDD D1 VSS VH VL SELD1 DVSS EF_AMUX21x
x3 VDD DVDD D2 VSS VH VL SELD2 DVSS EF_AMUX21x
x4 VDD DVDD D3 VSS VH VL SELD3 DVSS EF_AMUX21x
x5 VDD DVDD D4 VSS VH VL SELD4 DVSS EF_AMUX21x
x8 VDD DVDD D5 VSS VH VL SELD5 DVSS EF_AMUX21x
x9 VDD DVDD D6 VSS VH VL SELD6 DVSS EF_AMUX21x
x10 VDD DVDD D7 VSS VH VL SELD7 DVSS EF_AMUX21x
x11 VDD DVDD D8 VSS VH VL SELD8 DVSS EF_AMUX21x
x12 VDD DVDD D9 VSS VH VL SELD9 DVSS EF_AMUX21x
x6 VDD DVDD D10 VSS VH VL SELD10 DVSS EF_AMUX21x
x7 VDD DVDD D11 VSS VH VL SELD11 DVSS EF_AMUX21x
.ends


* expanding   symbol:  EF_SW_RST.sym # of pins=7
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SW_RST.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SW_RST.sch
.subckt EF_SW_RST VP1 VP2 AVDD DVDD AVSS RST DVSS
*.PININFO AVSS:B DVDD:B AVDD:B VP1:B VP2:B RST:I DVSS:B
x1 AVSS RST VP2 AVSS AVDD DVDD DVSS simple_analog_switch_ena1v8
x2 AVSS RST AVSS VP1 AVDD DVDD DVSS minimal_n_switch_ena1v8
.ends


* expanding   symbol:  EF_LSB_CAP.sym # of pins=8
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_LSB_CAP.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_LSB_CAP.sch
.subckt EF_LSB_CAP VP1 VSS D0 D1 D2 D3 D4 D5
*.PININFO VP1:B D0:B D1:B D2:B D3:B D4:B VSS:B D5:B
XC1 VP1 VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC2 VP1 D0 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=26
XC8 VSS VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VP1 D1 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC4 VP1 D2 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC5 VP1 D3 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC7 VP1 D4 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC9 D0 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC10 D1 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=2
XC11 D2 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XC12 D3 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=8
XC13 D4 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=16
XC14 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=26
XC15 VP1 D5 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC16 D5 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
.ends


* expanding   symbol:  EF_MSB_CAP.sym # of pins=8
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_MSB_CAP.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_MSB_CAP.sch
.subckt EF_MSB_CAP D8 D10 D9 VP2 D6 VSS D7 D11
*.PININFO D10:B D6:B D7:B D8:B D9:B VP2:B VSS:B D11:B
XC2 D6 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=27
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=27
XC6 VP2 D6 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC7 VP2 D7 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC8 VP2 D8 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC9 VP2 D9 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC10 VP2 D10 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC11 D7 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=2
XC12 D8 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XC13 D9 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=8
XC14 D10 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=16
XC1 VP2 D11 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC5 D11 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
.ends


* expanding   symbol:  EF_SC_CAP.sym # of pins=3
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SC_CAP.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_SC_CAP.sch
.subckt EF_SC_CAP VP1 VP2 VSS
*.PININFO VP1:B VP2:B VSS:B
XC13 VP1 VP2 sky130_fd_pr__cap_mim_m3_1 W=7 L=7.055 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7.055 m=9
XC1 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7.055 m=9
XC2 VP2 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7.055 m=1
.ends


* expanding   symbol:  EF_AMUX21x.sym # of pins=8
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX21x.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/xschem/EF_AMUX21x.sch
.subckt EF_AMUX21x vdd3p3 vdd1p8 vo vss a b sel dvss
*.PININFO sel:I vo:B vdd3p3:B vss:B vdd1p8:B dvss:B a:B b:B
x1 vss sel vo a vdd3p3 vdd1p8 dvss simple_analog_switch_ena1v8
x4 vss selp vo b vdd3p3 vdd1p8 dvss simple_analog_switch_ena1v8
x5 sel dvss dvss vdd1p8 vdd1p8 selp sky130_fd_sc_hd__inv_2
.ends


* expanding   symbol:  ../dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sym # of pins=7
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sch
.subckt simple_analog_switch_ena1v8 avss on out in avdd dvdd dvss
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B
x2 on dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
x3 net1 net2 avss out in avdd simple_analog_switch
x1 net3 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x4 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
x5[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  ../dependencies/sky130_ef_ip__analog_switches/xschem/minimal_n_switch_ena1v8.sym # of pins=7
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/minimal_n_switch_ena1v8.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/minimal_n_switch_ena1v8.sch
.subckt minimal_n_switch_ena1v8 avss on out in avdd dvdd dvss
*.PININFO on:I out:B in:B avdd:B dvdd:B dvss:B avss:B
x2 on dvdd dvss dvss avdd avdd net2 sky130_fd_sc_hvl__lsbuflv2hv_1
x1 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
x4 net1 dvss dvss avdd avdd net3 sky130_fd_sc_hvl__inv_2
x6 dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x3 net1 net3 out in avdd avss minimum_analog_switch
x5 on dvss dvss avdd avdd sky130_fd_sc_hvl__diode_2
.ends


* expanding   symbol:  simple_analog_switch.sym # of pins=6
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sch
.subckt simple_analog_switch on off vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B off:I
XM1 in on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 in off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=4 m=1
XM3 out off out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 out on out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM5 in off in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 in on in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
.ends


* expanding   symbol:  minimum_analog_switch.sym # of pins=6
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/minimum_analog_switch.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__cdac3v_12bit/dependencies/sky130_ef_ip__analog_switches/xschem/minimum_analog_switch.sch
.subckt minimum_analog_switch off on out in vdd vss
*.PININFO on:I out:B vss:B in:B off:I vdd:B
XM3 in off in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM1 out off out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=0.5 nf=1 m=1
XM4 out on in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=2 m=1
* noconn vdd
.ends

.end
