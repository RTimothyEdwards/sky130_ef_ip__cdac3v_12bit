magic
tech sky130A
magscale 1 2
timestamp 1717941056
<< metal3 >>
rect 85388 -19067 87868 -19003
rect 85388 -19191 87868 -19127
<< end >>
