magic
tech sky130A
magscale 1 2
timestamp 1718225130
<< error_s >>
rect 61184 11780 61265 11786
rect 61325 11780 61456 11786
rect 76064 11780 76145 11786
rect 76205 11780 76336 11786
rect 78544 11780 78625 11786
rect 78685 11780 78816 11786
rect 81024 11780 81105 11786
rect 81165 11780 81296 11786
rect 60944 11540 61184 11546
rect 61325 11540 61696 11546
rect 75824 11540 76064 11546
rect 76205 11540 76576 11546
rect 78304 11540 78544 11546
rect 78685 11540 79056 11546
rect 80784 11540 81024 11546
rect 81165 11540 81536 11546
rect 60894 11486 61265 11492
rect 61325 11486 61646 11492
rect 75774 11486 76145 11492
rect 76205 11486 76526 11492
rect 78254 11486 78625 11492
rect 78685 11486 79006 11492
rect 80734 11486 81105 11492
rect 81165 11486 81486 11492
rect 61134 11246 61265 11252
rect 61755 10843 61756 11389
rect 76014 11246 76145 11252
rect 76635 10843 76636 11389
rect 78494 11246 78625 11252
rect 79115 10843 79116 11389
rect 80974 11246 81105 11252
rect 81595 10843 81596 11389
rect 60425 10370 60485 10486
rect 62905 10370 62912 10486
rect 77785 10370 77845 10486
rect 80265 10370 80325 10486
rect 60027 10306 62912 10370
rect 75387 10306 82386 10370
rect 60027 10182 62912 10246
rect 75387 10182 82386 10246
rect 79465 10066 79525 10182
rect 60027 7826 60031 8197
rect 60079 7826 60085 8147
rect 60425 8015 60485 8130
rect 60417 7951 60493 8015
rect 60319 7890 60325 7907
rect 77785 7890 77845 8006
rect 82105 7890 82111 7957
rect 82345 7890 82351 8197
rect 60177 7826 60733 7890
rect 75387 7826 82386 7890
rect 60027 7445 60031 7766
rect 60079 7395 60085 7766
rect 60319 7635 60325 7766
rect 75387 7702 82386 7766
rect 76985 7586 77045 7702
rect 82105 7685 82111 7702
rect 79457 7577 79533 7641
rect 79465 7462 79525 7577
rect 81937 7576 82013 7640
rect 81942 7575 82008 7576
rect 81945 7462 82005 7575
rect 82345 7445 82351 7702
rect 81702 7335 82248 7336
rect 60027 5410 60031 5717
rect 60079 5410 60085 5667
rect 60425 5535 60485 5650
rect 60417 5471 60493 5535
rect 60319 5410 60325 5427
rect 62905 5410 62912 5526
rect 82105 5410 82111 5477
rect 82345 5410 82351 5717
rect 60027 5346 62912 5410
rect 75387 5346 82386 5410
rect 60027 5222 62912 5286
rect 75387 5222 82386 5286
rect 60027 4965 60031 5222
rect 60079 4915 60085 5222
rect 60319 5155 60325 5222
rect 79465 5106 79525 5222
rect 82105 5205 82111 5222
rect 81937 5096 82013 5160
rect 81942 5095 82008 5096
rect 81945 4982 82005 5095
rect 82345 4965 82351 5222
rect 81702 4855 82248 4856
rect 60027 2930 60031 3237
rect 60079 2930 60085 3187
rect 60425 3055 60485 3170
rect 60417 2991 60493 3055
rect 60319 2930 60325 2947
rect 62905 2930 62912 3046
rect 77785 2930 77845 3046
rect 82105 2930 82111 2997
rect 82345 2930 82351 3237
rect 60027 2866 62912 2930
rect 75387 2866 82386 2930
rect 60027 2742 62912 2806
rect 75387 2742 82386 2806
rect 60027 2485 60031 2742
rect 60079 2435 60085 2742
rect 60319 2675 60325 2742
rect 62105 2626 62165 2742
rect 79457 2617 79533 2681
rect 81945 2680 82005 2742
rect 82105 2725 82111 2742
rect 81937 2626 82013 2680
rect 79465 2502 79525 2617
rect 81937 2616 81945 2626
rect 82005 2616 82013 2626
rect 81942 2615 82008 2616
rect 82345 2485 82351 2742
rect 81702 2375 82248 2376
rect 60027 386 60031 757
rect 60079 386 60085 707
rect 60319 386 60325 467
rect 82105 440 82111 517
rect 81697 386 82253 440
rect 82345 386 82351 757
rect 60027 5 60031 326
rect 60079 -45 60085 326
rect 60319 195 60325 326
rect 82105 245 82111 326
rect 81937 146 82013 200
rect 81942 135 82008 136
rect 82345 5 82351 326
rect 81702 -105 82248 -104
rect 60027 -2094 60031 -1723
rect 60079 -2094 60085 -1773
rect 77785 -1905 77845 -1790
rect 60417 -1969 60493 -1914
rect 62897 -1969 62912 -1914
rect 77777 -1969 77853 -1905
rect 60319 -2094 60325 -2013
rect 80265 -2030 80325 -1914
rect 82105 -2030 82111 -1963
rect 82345 -2030 82351 -1723
rect 75387 -2094 82386 -2030
rect 60027 -2475 60031 -2154
rect 60079 -2525 60085 -2154
rect 60177 -2209 60733 -2154
rect 62657 -2209 62912 -2154
rect 60319 -2285 60325 -2209
rect 75387 -2218 82386 -2154
rect 79465 -2334 79525 -2218
rect 82105 -2235 82111 -2218
rect 81937 -2344 82013 -2280
rect 81942 -2345 82008 -2344
rect 81945 -2458 82005 -2345
rect 82345 -2475 82351 -2218
rect 81702 -2585 82248 -2584
rect 60027 -4574 60031 -4203
rect 60079 -4574 60085 -4253
rect 60425 -4385 60485 -4270
rect 60417 -4449 60493 -4385
rect 60319 -4510 60325 -4493
rect 77785 -4510 77845 -4394
rect 82105 -4510 82111 -4443
rect 82345 -4510 82351 -4203
rect 60177 -4574 60733 -4510
rect 75387 -4574 82386 -4510
rect 60027 -4955 60031 -4634
rect 60079 -5005 60085 -4634
rect 60319 -4765 60325 -4634
rect 75387 -4698 82386 -4634
rect 79465 -4814 79525 -4698
rect 82105 -4715 82111 -4698
rect 81937 -4824 82013 -4760
rect 81942 -4825 82008 -4824
rect 81945 -4938 82005 -4825
rect 82345 -4955 82351 -4698
rect 81702 -5065 82248 -5064
rect 60027 -6990 60031 -6683
rect 60079 -6990 60085 -6733
rect 60425 -6865 60485 -6750
rect 62905 -6865 62912 -6750
rect 77785 -6865 77845 -6750
rect 60417 -6929 60493 -6865
rect 62897 -6929 62912 -6865
rect 77777 -6929 77853 -6865
rect 60319 -6990 60325 -6973
rect 82105 -6990 82111 -6923
rect 82345 -6990 82351 -6683
rect 60027 -7054 62912 -6990
rect 75387 -7054 82386 -6990
rect 60027 -7178 62912 -7114
rect 75387 -7178 82386 -7114
rect 60027 -7435 60031 -7178
rect 60079 -7485 60085 -7178
rect 60319 -7245 60325 -7178
rect 79465 -7294 79525 -7178
rect 82105 -7195 82111 -7178
rect 81937 -7304 82013 -7240
rect 81942 -7305 82008 -7304
rect 81945 -7418 82005 -7305
rect 82345 -7435 82351 -7178
rect 81702 -7545 82248 -7544
rect 60027 -9534 60031 -9163
rect 60079 -9534 60085 -9213
rect 60425 -9345 60485 -9230
rect 60417 -9409 60493 -9345
rect 60319 -9470 60325 -9453
rect 60177 -9534 60733 -9470
rect 82105 -9480 82111 -9403
rect 81697 -9534 82253 -9480
rect 82345 -9534 82351 -9163
rect 60027 -9915 60031 -9594
rect 60079 -9965 60085 -9594
rect 60319 -9725 60325 -9594
rect 82105 -9675 82111 -9594
rect 81937 -9774 82013 -9720
rect 81942 -9785 82008 -9784
rect 82345 -9915 82351 -9594
rect 81702 -10025 82248 -10024
rect 61263 -10310 61327 -10268
rect 76143 -10310 76207 -10268
rect 78623 -10310 78687 -10268
rect 81103 -10310 81167 -10268
rect 61184 -10496 61263 -10310
rect 61327 -10496 61456 -10310
rect 76064 -10496 76143 -10310
rect 76207 -10496 76336 -10310
rect 78544 -10496 78623 -10310
rect 78687 -10496 78816 -10310
rect 81024 -10496 81103 -10310
rect 81167 -10496 81296 -10310
rect 61263 -10540 61327 -10496
rect 76143 -10540 76207 -10496
rect 78623 -10540 78687 -10496
rect 81103 -10540 81167 -10496
rect 61265 -10550 61325 -10540
rect 76145 -10550 76205 -10540
rect 78625 -10550 78685 -10540
rect 81105 -10550 81165 -10540
rect 61265 -11090 61325 -11077
rect 76145 -11090 76205 -11077
rect 78625 -11090 78685 -11077
rect 81105 -11090 81165 -11077
rect 61263 -11131 61327 -11090
rect 76143 -11131 76207 -11090
rect 78623 -11131 78687 -11090
rect 81103 -11131 81167 -11090
rect 61134 -11317 61263 -11131
rect 61327 -11317 61406 -11131
rect 76014 -11317 76143 -11131
rect 76207 -11317 76286 -11131
rect 78494 -11317 78623 -11131
rect 78687 -11317 78766 -11131
rect 80974 -11317 81103 -11131
rect 81167 -11317 81246 -11131
rect 61263 -11362 61327 -11317
rect 76143 -11362 76207 -11317
rect 78623 -11362 78687 -11317
rect 81103 -11362 81167 -11317
rect 60182 -11606 60728 -11605
rect 60027 -12036 60031 -11665
rect 60079 -12036 60085 -11715
rect 60422 -11846 60488 -11845
rect 60417 -11910 60493 -11856
rect 60319 -12036 60325 -11955
rect 82105 -12036 82111 -11905
rect 82345 -12036 82351 -11665
rect 60027 -12417 60031 -12096
rect 60079 -12467 60085 -12096
rect 60177 -12150 60733 -12096
rect 60319 -12227 60325 -12150
rect 81697 -12160 82253 -12096
rect 82105 -12177 82111 -12160
rect 81937 -12286 82013 -12222
rect 81942 -12287 82008 -12286
rect 81945 -12400 82005 -12287
rect 82345 -12417 82351 -12096
rect 81702 -12527 82248 -12526
rect 77785 -14452 77845 -14336
rect 82105 -14452 82111 -14385
rect 82345 -14452 82351 -14145
rect 75387 -14516 82386 -14452
rect 75387 -14640 82386 -14576
rect 76985 -14756 77045 -14640
rect 82105 -14657 82111 -14640
rect 79457 -14765 79533 -14701
rect 79465 -14880 79525 -14765
rect 81937 -14766 82013 -14702
rect 81942 -14767 82008 -14766
rect 81945 -14880 82005 -14767
rect 82345 -14897 82351 -14640
rect 81702 -15007 82248 -15006
rect 75387 -16996 77042 -16932
rect 82105 -16996 82111 -16865
rect 82345 -16996 82351 -16625
rect 75387 -17120 77042 -17056
rect 81697 -17120 82253 -17056
rect 82105 -17137 82111 -17120
rect 81937 -17246 82013 -17182
rect 81942 -17247 82008 -17246
rect 81945 -17360 82005 -17247
rect 82345 -17377 82351 -17056
rect 81702 -17487 82248 -17486
rect 79217 -19476 79773 -19421
rect 82105 -19422 82111 -19345
rect 81697 -19476 82253 -19422
rect 82345 -19476 82351 -19105
rect 82105 -19617 82111 -19536
rect 79457 -19716 79533 -19661
rect 81937 -19716 82013 -19662
rect 81942 -19727 82008 -19726
rect 82345 -19857 82351 -19536
rect 81702 -19967 82248 -19966
rect 77777 -21831 77853 -21776
rect 75387 -21956 77042 -21892
rect 82105 -21956 82111 -21825
rect 82345 -21956 82351 -21585
rect 75387 -22080 77042 -22016
rect 77537 -22071 78093 -22016
rect 81697 -22080 82253 -22016
rect 82105 -22097 82111 -22080
rect 81937 -22206 82013 -22142
rect 81942 -22207 82008 -22206
rect 81945 -22320 82005 -22207
rect 82345 -22337 82351 -22016
rect 81702 -22447 82248 -22446
rect 77785 -24247 77845 -24132
rect 77777 -24311 77853 -24247
rect 80265 -24372 80325 -24256
rect 82105 -24372 82111 -24305
rect 82345 -24372 82351 -24065
rect 75387 -24436 82386 -24372
rect 75387 -24560 82386 -24496
rect 79465 -24676 79525 -24560
rect 82105 -24577 82111 -24560
rect 81937 -24686 82013 -24622
rect 81942 -24687 82008 -24686
rect 81945 -24800 82005 -24687
rect 82345 -24817 82351 -24560
rect 81702 -24927 82248 -24926
rect 77785 -26852 77845 -26736
rect 82105 -26852 82111 -26785
rect 82345 -26852 82351 -26545
rect 75387 -26916 82386 -26852
rect 75387 -27040 82386 -26976
rect 79465 -27156 79525 -27040
rect 82105 -27057 82111 -27040
rect 81937 -27166 82013 -27102
rect 81942 -27167 82008 -27166
rect 81945 -27280 82005 -27167
rect 82345 -27297 82351 -27040
rect 81702 -27407 82248 -27406
rect 77785 -29207 77845 -29092
rect 77777 -29271 77853 -29207
rect 82105 -29332 82111 -29265
rect 82345 -29332 82351 -29025
rect 75387 -29396 82386 -29332
rect 75387 -29520 82386 -29456
rect 60027 -29777 60031 -29626
rect 60079 -29827 60085 -29626
rect 79465 -29636 79525 -29520
rect 82105 -29537 82111 -29520
rect 81937 -29646 82013 -29582
rect 81942 -29647 82008 -29646
rect 81945 -29760 82005 -29647
rect 82345 -29777 82351 -29520
rect 81702 -29887 82248 -29886
rect 62905 -31812 62912 -31696
rect 77785 -31812 77845 -31696
rect 60027 -31876 62912 -31812
rect 75387 -31876 82386 -31812
rect 60027 -32000 62912 -31936
rect 75387 -32000 82386 -31936
rect 62105 -32116 62165 -32000
rect 76985 -32116 77045 -32000
rect 79465 -32116 79525 -32000
rect 81945 -32116 82005 -32000
rect 61184 -32882 61265 -32876
rect 61325 -32882 61456 -32876
rect 76064 -32882 76145 -32876
rect 76205 -32882 76336 -32876
rect 78544 -32882 78625 -32876
rect 78685 -32882 78816 -32876
rect 81024 -32882 81105 -32876
rect 81165 -32882 81296 -32876
rect 60944 -33122 61184 -33116
rect 61325 -33122 61696 -33116
rect 75824 -33122 76064 -33116
rect 76205 -33122 76576 -33116
rect 78304 -33122 78544 -33116
rect 78685 -33122 79056 -33116
rect 80784 -33122 81024 -33116
rect 81165 -33122 81536 -33116
rect 60894 -33176 61265 -33170
rect 61325 -33176 61646 -33170
rect 75774 -33176 76145 -33170
rect 76205 -33176 76526 -33170
rect 78254 -33176 78625 -33170
rect 78685 -33176 79006 -33170
rect 80734 -33176 81105 -33170
rect 81165 -33176 81486 -33170
rect 61134 -33416 61265 -33410
rect 61755 -33819 61756 -33273
rect 76014 -33416 76145 -33410
rect 76635 -33819 76636 -33273
rect 78494 -33416 78625 -33410
rect 79115 -33819 79116 -33273
rect 80974 -33416 81105 -33410
rect 81595 -33819 81596 -33273
<< viali >>
rect 58720 12899 83690 12933
rect 58631 -34472 58665 12845
rect 83747 -34470 83781 12837
rect 58722 -34559 83692 -34525
<< metal1 >>
rect 53524 14365 68765 14413
rect 53335 14269 70877 14317
rect 71172 14269 89082 14317
rect 53239 14173 69361 14221
rect 69662 14173 89177 14221
rect 53142 14077 70117 14125
rect 70415 14077 89273 14125
rect 53046 13981 72767 14029
rect 76033 13981 89368 14029
rect 76033 13933 76081 13981
rect 52949 13885 68727 13933
rect 72328 13885 76081 13933
rect 76152 13885 89464 13933
rect 68679 13837 68727 13885
rect 52849 13789 68605 13837
rect 68679 13789 72007 13837
rect 68557 13645 68605 13789
rect 76152 13741 76200 13885
rect 71570 13693 76200 13741
rect 76267 13789 89562 13837
rect 68557 13597 73528 13645
rect 76267 13549 76315 13789
rect 73085 13501 76315 13549
rect 58611 12933 83801 12953
rect 58611 12899 58720 12933
rect 83690 12899 83801 12933
rect 58611 12879 83801 12899
rect 58611 12845 58685 12879
rect 52856 8734 53526 8782
rect 52952 1730 53526 1778
rect 53048 -5275 53526 -5227
rect 53089 -19283 53526 -19235
rect 53089 -26286 53526 -26238
rect 53089 -33290 53526 -33242
rect 58611 -34472 58631 12845
rect 58665 -34472 58685 12845
rect 58611 -34505 58685 -34472
rect 83727 12837 83801 12879
rect 83727 -34470 83747 12837
rect 83781 -34470 83801 12837
rect 88887 8733 89557 8781
rect 88887 1730 89469 1778
rect 88887 -5274 89372 -5226
rect 88887 -19282 89306 -19234
rect 88886 -26286 89322 -26238
rect 88887 -33290 89322 -33242
rect 83727 -34505 83801 -34470
rect 58611 -34525 83801 -34505
rect 58611 -34559 58722 -34525
rect 83692 -34559 83801 -34525
rect 58611 -34579 83801 -34559
rect 58611 -34690 58685 -34579
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -34948 58685 -34939
rect 83727 -34698 83801 -34579
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 83727 -34955 83801 -34947
<< via1 >>
rect 58619 -34939 58678 -34690
rect 83734 -34947 83793 -34698
<< metal2 >>
rect 53488 14421 53565 14432
rect 52859 8730 52907 13786
rect 52955 1725 53003 13940
rect 53051 -5279 53099 14037
rect 53147 -19329 53195 14131
rect 53243 -26299 53291 14225
rect 53339 -33302 53387 14325
rect 53488 14235 53498 14421
rect 53555 14235 53565 14421
rect 53488 14224 53565 14235
rect 67192 13923 68325 14589
rect 68837 14413 69037 14589
rect 68765 14365 69037 14413
rect 69217 14389 69417 14589
rect 69602 14390 69802 14590
rect 69980 14391 70180 14591
rect 70363 14391 70563 14591
rect 70742 14391 70942 14591
rect 69294 14158 69342 14389
rect 69674 14158 69722 14390
rect 70054 14067 70102 14391
rect 70434 14067 70482 14391
rect 70814 14259 70862 14391
rect 71124 14389 71324 14589
rect 71501 14391 71701 14591
rect 71886 14391 72086 14591
rect 72256 14391 72456 14591
rect 72639 14391 72839 14591
rect 71194 14259 71242 14389
rect 67192 13577 67221 13923
rect 68290 13577 68325 13923
rect 71574 13692 71622 14391
rect 71954 13788 72002 14391
rect 72334 13881 72382 14391
rect 72714 13975 72762 14391
rect 73014 14389 73214 14589
rect 73392 14391 73592 14591
rect 74028 14498 75160 14592
rect 67192 13552 68325 13577
rect 73094 13494 73142 14389
rect 73474 13588 73522 14391
rect 74028 14149 74053 14498
rect 75137 14149 75160 14498
rect 74028 14123 75160 14149
rect 57639 -9376 57703 -7904
rect 53490 -9387 53561 -9377
rect 53490 -9561 53498 -9387
rect 53555 -9561 53561 -9387
rect 53490 -9570 53561 -9561
rect 57639 -9667 57703 -9658
rect 57639 -11972 57703 -11963
rect 57639 -13726 57703 -12254
rect 89029 -33326 89077 14327
rect 89125 -26323 89173 14226
rect 89221 -19307 89269 14132
rect 89317 -5309 89365 14033
rect 89413 1725 89461 13938
rect 89509 8726 89557 13844
rect 58611 -34690 58685 -34682
rect 58611 -34939 58619 -34690
rect 58678 -34939 58685 -34690
rect 58611 -36347 58685 -34939
rect 83727 -34698 83801 -34690
rect 83727 -34947 83734 -34698
rect 83793 -34947 83801 -34698
rect 68751 -35760 70341 -35717
rect 68751 -36098 68783 -35760
rect 70303 -36098 70341 -35760
rect 58611 -36358 58735 -36347
rect 58611 -36734 58624 -36358
rect 58724 -36734 58735 -36358
rect 58611 -36741 58735 -36734
rect 58612 -36746 58735 -36741
rect 68751 -36856 70341 -36098
rect 72201 -36381 73791 -36342
rect 83727 -36347 83801 -34947
rect 72201 -36719 72237 -36381
rect 73757 -36719 73791 -36381
rect 72201 -36868 73791 -36719
rect 83672 -36359 83801 -36347
rect 83672 -36735 83686 -36359
rect 83789 -36735 83801 -36359
rect 83672 -36747 83801 -36735
<< via2 >>
rect 53498 14235 53555 14421
rect 67221 13577 68290 13923
rect 74053 14149 75137 14498
rect 53498 -9561 53555 -9387
rect 57639 -9658 57703 -9376
rect 57639 -12254 57703 -11972
rect 68783 -36098 70303 -35760
rect 58624 -36734 58724 -36358
rect 72237 -36719 73757 -36381
rect 83686 -36735 83789 -36359
<< metal3 >>
rect 53488 14421 53565 14432
rect 53488 14235 53498 14421
rect 53555 14235 53565 14421
rect 53488 14224 53565 14235
rect 53496 -9377 53556 14224
rect 65040 14202 65240 14402
rect 64616 13678 64816 13878
rect 57444 10306 57452 10370
rect 57681 10306 58425 10370
rect 84059 10182 85236 10246
rect 57196 7826 58405 7890
rect 57189 2742 58413 2806
rect 83551 2742 84399 2806
rect 84606 2742 84613 2806
rect 83933 262 85241 326
rect 57199 -4698 58320 -4634
rect 85203 -6990 85398 -6851
rect 83918 -7054 85398 -6990
rect 57634 -9376 57708 -9370
rect 53490 -9387 53561 -9377
rect 53490 -9561 53498 -9387
rect 53555 -9561 53561 -9387
rect 53490 -9570 53561 -9561
rect 57634 -9658 57639 -9376
rect 57703 -9594 57708 -9376
rect 88726 -9586 88955 -9580
rect 85166 -9594 85373 -9588
rect 57703 -9658 58900 -9594
rect 83980 -9658 85171 -9594
rect 85367 -9658 85373 -9594
rect 57634 -9663 57708 -9658
rect 85166 -9664 85373 -9658
rect 88726 -9661 88735 -9586
rect 88946 -9594 88955 -9586
rect 89380 -9594 89580 -9508
rect 88946 -9658 89580 -9594
rect 88946 -9661 88955 -9658
rect 88726 -9668 88955 -9661
rect 89380 -9708 89580 -9658
rect 88726 -11966 88955 -11960
rect 57634 -11972 57708 -11967
rect 85166 -11972 85372 -11967
rect 57634 -12254 57639 -11972
rect 57703 -12036 58919 -11972
rect 83980 -12036 85170 -11972
rect 85366 -12036 85372 -11972
rect 57703 -12254 57708 -12036
rect 85166 -12041 85372 -12036
rect 88726 -12041 88736 -11966
rect 88947 -11972 88955 -11966
rect 89380 -11972 89577 -11889
rect 88947 -12036 89577 -11972
rect 88947 -12041 88955 -12036
rect 88726 -12048 88955 -12041
rect 89380 -12089 89577 -12036
rect 57634 -12260 57708 -12254
rect 57014 -14640 58370 -14576
rect 57014 -14663 57210 -14640
rect 83950 -16996 85256 -16932
rect 57162 -21956 58447 -21892
rect 54633 -24342 55033 -24324
rect 54633 -24464 54649 -24342
rect 55017 -24464 55033 -24342
rect 58042 -24368 58280 -24356
rect 58042 -24434 58054 -24368
rect 58266 -24372 58280 -24368
rect 58266 -24434 58410 -24372
rect 58042 -24436 58410 -24434
rect 83988 -24436 85241 -24372
rect 58042 -24450 58280 -24436
rect 54633 -24480 55033 -24464
rect 83963 -29520 85239 -29456
rect 57194 -31876 58330 -31812
rect 83980 -32000 84409 -31936
rect 84644 -32000 84651 -31936
rect 70647 -35210 70847 -35010
rect 71047 -35490 71247 -35290
rect 65838 -36033 66038 -35833
rect 65303 -36648 65503 -36448
<< via3 >>
rect 54639 10282 55027 10405
rect 57452 10306 57681 10370
rect 84399 2742 84606 2806
rect 87392 2709 87769 2840
rect 85171 -9658 85367 -9594
rect 88735 -9661 88946 -9586
rect 85170 -12036 85366 -11972
rect 88736 -12041 88947 -11966
rect 54649 -24464 55017 -24342
rect 58054 -24434 58266 -24368
rect 84409 -32000 84644 -31936
rect 87386 -32019 87774 -31915
<< metal4 >>
rect 54633 10405 55033 10406
rect 54633 10282 54639 10405
rect 55027 10370 55033 10405
rect 57451 10370 57682 10371
rect 55027 10306 57452 10370
rect 57681 10306 57682 10370
rect 55027 10282 55033 10306
rect 57451 10305 57682 10306
rect 54633 10281 55033 10282
rect 87380 2840 87780 2851
rect 84398 2806 84607 2807
rect 87380 2806 87392 2840
rect 84398 2742 84399 2806
rect 84606 2742 87392 2806
rect 84398 2741 84607 2742
rect 87380 2709 87392 2742
rect 87769 2709 87780 2840
rect 87380 2697 87780 2709
rect 88726 -9586 88955 -9580
rect 85166 -9594 85373 -9588
rect 88726 -9594 88735 -9586
rect 85166 -9658 85171 -9594
rect 85367 -9658 88735 -9594
rect 85166 -9664 85373 -9658
rect 88726 -9661 88735 -9658
rect 88946 -9661 88955 -9586
rect 88726 -9668 88955 -9661
rect 88726 -11966 88955 -11960
rect 85166 -11972 85372 -11967
rect 88726 -11972 88736 -11966
rect 85166 -12036 85170 -11972
rect 85366 -12036 88736 -11972
rect 85166 -12041 85372 -12036
rect 88726 -12041 88736 -12036
rect 88947 -12041 88955 -11966
rect 88726 -12048 88955 -12041
rect 54631 -24342 55037 -24324
rect 54631 -24464 54649 -24342
rect 55017 -24374 55037 -24342
rect 58042 -24368 58280 -24356
rect 58042 -24374 58054 -24368
rect 55017 -24434 58054 -24374
rect 58266 -24434 58280 -24368
rect 55017 -24464 55037 -24434
rect 58042 -24450 58280 -24434
rect 54631 -24480 55037 -24464
rect 87380 -31915 87780 -31914
rect 84408 -31936 84645 -31935
rect 87380 -31936 87386 -31915
rect 84408 -32000 84409 -31936
rect 84644 -32000 87386 -31936
rect 84408 -32001 84645 -32000
rect 87380 -32019 87386 -32000
rect 87774 -32019 87780 -31915
rect 87380 -32020 87780 -32019
use cdac_dummy_switch  cdac_dummy_switch_1
timestamp 1718223925
transform -1 0 133337 0 1 6988
box 44011 -15952 48431 -14149
use cdac_dummy_switch  cdac_dummy_switch_2
timestamp 1718223925
transform -1 0 133337 0 -1 -28520
box 44011 -15952 48431 -14149
use cdac_via_3cut  cdac_via_3cut_0
timestamp 1718157421
transform 1 0 212 0 1 34864
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_1
timestamp 1718157421
transform 1 0 597 0 1 -156
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_2
timestamp 1718157421
transform 1 0 501 0 1 6844
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_3
timestamp 1718157421
transform 1 0 405 0 1 13803
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_4
timestamp 1718157421
transform 1 0 308 0 1 27859
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_5
timestamp 1718157421
transform 1 0 36481 0 1 13852
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_6
timestamp 1718157421
transform 1 0 116 0 1 41869
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_7
timestamp 1718157421
transform 1 0 36286 0 1 -156
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_8
timestamp 1718157421
transform 1 0 36382 0 1 6846
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_9
timestamp 1718157421
transform 1 0 36571 0 1 27862
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_10
timestamp 1718157421
transform 1 0 36767 0 1 41869
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_11
timestamp 1718157421
transform 1 0 36670 0 1 34866
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_12
timestamp 1718157421
transform 1 0 116 0 1 46924
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_13
timestamp 1718157421
transform 1 0 213 0 1 47021
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_14
timestamp 1718157421
transform 1 0 308 0 1 47117
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_15
timestamp 1718157421
transform 1 0 404 0 1 47213
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_16
timestamp 1718157421
transform 1 0 501 0 1 47308
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_17
timestamp 1718157421
transform 1 0 595 0 1 47403
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_18
timestamp 1718157421
transform 1 0 36768 0 1 46925
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_19
timestamp 1718157421
transform 1 0 36670 0 1 47019
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_20
timestamp 1718157421
transform 1 0 36574 0 1 47117
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_21
timestamp 1718157421
transform 1 0 36478 0 1 47212
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_22
timestamp 1718157421
transform 1 0 36381 0 1 47309
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_23
timestamp 1718157421
transform 1 0 36286 0 1 47405
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_24
timestamp 1718157421
transform 0 1 103797 -1 0 67058
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_25
timestamp 1718157421
transform 0 1 102275 -1 0 66961
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_26
timestamp 1718157421
transform 0 1 104329 -1 0 67057
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_27
timestamp 1718157421
transform 0 1 103040 -1 0 66865
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_28
timestamp 1718157421
transform 0 1 102807 -1 0 66959
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_29
timestamp 1718157421
transform 0 1 103566 -1 0 66867
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_30
timestamp 1718157421
transform 0 1 104707 -1 0 66480
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_31
timestamp 1718157421
transform 0 1 105697 -1 0 66770
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_32
timestamp 1718157421
transform 0 1 105466 -1 0 66677
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_33
timestamp 1718157421
transform 0 1 104940 -1 0 66579
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_34
timestamp 1718157421
transform 0 1 106228 -1 0 66291
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_35
timestamp 1718157421
transform 0 1 106453 -1 0 66386
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_36
timestamp 1718157421
transform 0 1 86645 -1 0 67155
box 52740 -33138 52792 -32927
use cdac_via_3cut  cdac_via_3cut_37
timestamp 1718157421
transform 0 1 101701 -1 0 67154
box 52740 -33138 52792 -32927
use EF_SW_RST  x1
timestamp 1718225130
transform 1 0 52769 0 -1 -10037
box 250 -2876 4934 4334
use EF_AMUX0201_ARRAY1  x3
timestamp 1718225130
transform 0 1 62083 -1 0 14841
box 320 -9064 51588 27311
use EF_BANK_CAP_12  x4
timestamp 1718225130
transform 1 0 0 0 1 -8000
box 58243 -26645 84124 21019
<< labels >>
flabel metal3 64616 13678 64816 13878 0 FreeSans 256 90 0 0 DVSS
port 12 nsew
flabel metal3 71047 -35490 71247 -35290 0 FreeSans 256 90 0 0 VH
port 14 nsew
flabel metal3 70647 -35210 70847 -35010 0 FreeSans 256 90 0 0 VL
port 15 nsew
flabel metal3 65838 -36033 66038 -35833 0 FreeSans 256 90 0 0 VSS
port 13 nsew
flabel metal3 65303 -36648 65503 -36448 0 FreeSans 256 90 0 0 VDD
port 10 nsew
flabel metal3 65040 14202 65240 14402 0 FreeSans 256 90 0 0 DVDD
port 11 nsew
flabel metal3 89380 -9708 89580 -9508 0 FreeSans 480 0 0 0 OUT
port 16 nsew
flabel metal3 89380 -12089 89577 -11889 0 FreeSans 480 0 0 0 OUTNC
port 22 nsew
flabel metal2 71501 14391 71701 14591 0 FreeSans 480 0 0 0 SELD6
port 6 nsew
flabel metal2 73392 14391 73592 14591 0 FreeSans 480 0 0 0 SELD11
port 21 nsew
flabel metal2 73014 14389 73214 14589 0 FreeSans 480 0 0 0 SELD10
port 19 nsew
flabel metal2 72639 14391 72839 14591 0 FreeSans 480 0 0 0 SELD9
port 9 nsew
flabel metal2 71886 14391 72086 14591 0 FreeSans 480 0 0 0 SELD7
port 7 nsew
flabel metal2 72256 14391 72456 14591 0 FreeSans 480 0 0 0 SELD8
port 8 nsew
flabel metal2 69980 14391 70180 14591 0 FreeSans 480 0 0 0 SELD2
port 2 nsew
flabel metal2 70363 14391 70563 14591 0 FreeSans 480 0 0 0 SELD3
port 3 nsew
flabel metal2 70742 14391 70942 14591 0 FreeSans 480 0 0 0 SELD4
port 4 nsew
flabel metal2 71124 14389 71324 14589 0 FreeSans 480 0 0 0 SELD5
port 5 nsew
flabel metal2 69602 14390 69802 14590 0 FreeSans 480 0 0 0 SELD1
port 24 nsew
flabel metal2 69217 14389 69417 14589 0 FreeSans 480 0 0 0 SELD0
port 23 nsew
flabel metal2 68837 14389 69037 14589 0 FreeSans 480 0 0 0 RST
port 17 nsew
<< end >>
