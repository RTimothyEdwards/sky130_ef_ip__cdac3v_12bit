magic
tech sky130A
magscale 1 2
timestamp 1718247631
<< error_p >>
rect 83248 -26401 83568 -26353
rect 83248 -26637 83290 -26401
rect 83248 -26673 83568 -26637
<< metal3 >>
rect 84178 -26318 84238 -26177
rect 84170 -26382 84176 -26318
rect 84240 -26382 84246 -26318
rect 82568 -26507 85050 -26443
rect 82568 -26631 83291 -26567
rect 83525 -26631 84176 -26567
rect 84240 -26631 85050 -26567
<< via3 >>
rect 84176 -26382 84240 -26318
rect 83291 -26631 83525 -26567
rect 84176 -26631 84240 -26567
<< metal4 >>
rect 84174 -26318 84241 -26317
rect 84174 -26382 84176 -26318
rect 84240 -26382 84241 -26318
rect 84174 -26567 84241 -26382
rect 84174 -26631 84176 -26567
rect 84240 -26631 84241 -26567
rect 84174 -26632 84241 -26631
<< via4 >>
rect 83290 -26567 83526 -26401
rect 83290 -26631 83291 -26567
rect 83291 -26631 83525 -26567
rect 83525 -26631 83526 -26567
rect 83290 -26637 83526 -26631
<< metal5 >>
rect 83248 -26401 83568 -26362
rect 83248 -26637 83290 -26401
rect 83526 -26637 83568 -26401
rect 83248 -26673 83568 -26637
<< end >>
