magic
tech sky130A
magscale 1 2
timestamp 1718157421
<< checkpaint >>
rect 52740 -33138 52792 -32927
<< metal1 >>
rect 52740 -32934 52792 -32927
rect 52740 -33138 52792 -33131
<< via1 >>
rect 52740 -33131 52792 -32934
<< metal2 >>
rect 52740 -32934 52792 -32927
rect 52740 -33138 52792 -33131
<< end >>
