magic
tech sky130A
magscale 1 2
timestamp 1717948824
<< metal1 >>
rect 83461 -2699 83661 -2499
rect 58660 -3406 58860 -3206
rect 58666 -13946 58866 -13746
rect 58614 -16437 58814 -16237
rect 58092 -17622 58292 -17422
rect 58092 -18422 58292 -18222
rect 58092 -19222 58292 -19022
rect 58092 -19622 58292 -19422
rect 58092 -20022 58292 -19822
rect 58092 -20822 58292 -20622
rect 58092 -21222 58292 -21022
rect 58092 -22022 58292 -21822
rect 58092 -22422 58292 -22222
<< via3 >>
rect 72347 10742 72565 10806
rect 69860 -1658 70081 -1594
<< metal4 >>
rect 72346 10806 72566 10807
rect 72346 10742 72347 10806
rect 72565 10742 72566 10806
rect 72346 10741 72566 10742
rect 72425 10476 72485 10741
rect 60025 -1924 60085 -1204
rect 69945 -1593 70005 -1144
rect 69859 -1594 70082 -1593
rect 69859 -1658 69860 -1594
rect 70081 -1658 70082 -1594
rect 69859 -1659 70082 -1658
rect 82345 -1924 82405 -1204
rect 60935 -2845 61655 -2785
rect 63415 -2845 64135 -2785
rect 65895 -2845 66615 -2785
rect 73335 -2845 74055 -2785
rect 75815 -2845 76535 -2785
rect 78295 -2845 79015 -2785
rect 80775 -2845 81495 -2785
rect 60025 -4426 60085 -3706
rect 69945 -4426 70005 -3705
rect 82345 -4426 82405 -3706
rect 69945 -14346 70005 -13626
rect 68375 -15256 69095 -15196
rect 70855 -15256 71575 -15196
rect 69945 -16826 70005 -16106
use cap_array_half  cap_array_half_0
timestamp 1717946239
transform -1 0 164043 0 -1 -5781
box 80293 -26673 105363 -4081
use cap_array_half  cap_array_half_1
timestamp 1717946239
transform 1 0 -21613 0 1 151
box 80293 -26673 105363 -4081
use caparray_connect_near  caparray_connect_near_0
timestamp 1717937330
transform -1 0 151643 0 -1 -28101
box 80427 -26673 82908 -26177
use cdac_ratioed_cap  cdac_ratioed_cap_0
array 0 9 2480 0 0 2797
timestamp 1717944067
transform 1 0 -21716 0 1 29649
box 80396 -33851 83146 -31078
<< labels >>
flabel metal1 58092 -17622 58292 -17422 0 FreeSans 256 0 0 0 D8
port 0 nsew
flabel metal1 58092 -18422 58292 -18222 0 FreeSans 256 0 0 0 D4
port 2 nsew
flabel metal1 58092 -19222 58292 -19022 0 FreeSans 256 0 0 0 D9
port 4 nsew
flabel metal1 58092 -19622 58292 -19422 0 FreeSans 256 0 0 0 D5
port 5 nsew
flabel metal1 58092 -20022 58292 -19822 0 FreeSans 256 0 0 0 D1
port 6 nsew
flabel metal1 58092 -20822 58292 -20622 0 FreeSans 256 0 0 0 D2
port 8 nsew
flabel metal1 58092 -21222 58292 -21022 0 FreeSans 256 0 0 0 D6
port 9 nsew
flabel metal1 58092 -22022 58292 -21822 0 FreeSans 256 0 0 0 D7
port 11 nsew
flabel metal1 58092 -22422 58292 -22222 0 FreeSans 256 0 0 0 D3
port 12 nsew
flabel metal1 58614 -16437 58814 -16237 0 FreeSans 256 0 0 0 VSS
port 10 nsew
flabel metal1 58666 -13946 58866 -13746 0 FreeSans 256 0 0 0 D0
port 1 nsew
flabel metal1 58660 -3406 58860 -3206 0 FreeSans 256 0 0 0 VP1
port 3 nsew
flabel metal1 83461 -2699 83661 -2499 0 FreeSans 256 0 0 0 VP2
port 7 nsew
<< end >>
