magic
tech sky130A
magscale 1 2
timestamp 1718210529
<< dnwell >>
rect 58654 -26536 83758 20910
<< nwell >>
rect 58545 20704 83867 21019
rect 58545 -26330 58860 20704
rect 83552 -26330 83867 20704
rect 58545 -26645 83867 -26330
<< mvnsubdiff >>
rect 58611 20933 83801 20953
rect 58611 20899 58691 20933
rect 83721 20899 83801 20933
rect 58611 20879 83801 20899
rect 58611 20873 58685 20879
rect 58611 -26499 58631 20873
rect 58665 -26499 58685 20873
rect 58611 -26505 58685 -26499
rect 83727 20873 83801 20879
rect 83727 -26499 83747 20873
rect 83781 -26499 83801 20873
rect 83727 -26505 83801 -26499
rect 58611 -26525 83801 -26505
rect 58611 -26559 58691 -26525
rect 83721 -26559 83801 -26525
rect 58611 -26579 83801 -26559
<< mvnsubdiffcont >>
rect 58691 20899 83721 20933
rect 58631 -26499 58665 20873
rect 83747 -26499 83781 20873
rect 58691 -26559 83721 -26525
<< locali >>
rect 58611 20933 83801 20953
rect 58611 20899 58691 20933
rect 83721 20899 83801 20933
rect 58611 20879 83801 20899
rect 58611 20873 58685 20879
rect 58611 -26499 58631 20873
rect 58665 -26499 58685 20873
rect 58611 -26505 58685 -26499
rect 83727 20873 83801 20879
rect 83727 -26499 83747 20873
rect 83781 -26499 83801 20873
rect 83727 -26505 83801 -26499
rect 58611 -26525 83801 -26505
rect 58611 -26559 58691 -26525
rect 83721 -26559 83801 -26525
rect 58611 -26579 83801 -26559
<< metal3 >>
rect 58361 18306 58817 18370
rect 83378 18182 83379 18246
rect 83445 18182 83446 18246
rect 83523 18182 84124 18246
rect 58323 15826 58917 15890
rect 58987 15826 58988 15890
rect 59052 15826 59053 15890
rect 83503 15702 83504 15766
rect 83568 15702 83569 15766
rect 58865 13346 58866 13410
rect 58930 13346 58931 13410
rect 83378 13222 83379 13286
rect 83445 13222 83446 13286
rect 58988 10866 58989 10930
rect 59053 10866 59054 10930
rect 58342 10742 58743 10806
rect 58807 10742 58980 10806
rect 81945 10552 82005 10776
rect 58865 8386 58866 8450
rect 58930 8386 58931 8450
rect 83445 8262 83997 8326
rect 58737 5906 58743 5970
rect 58807 5906 58879 5970
rect 58988 5782 58989 5846
rect 59053 5782 59054 5846
rect 83378 3426 83379 3490
rect 83445 3426 83446 3490
rect 58256 3302 58866 3366
rect 58930 3302 59007 3366
rect 83448 946 83504 1010
rect 83568 946 83982 1010
rect 83534 -1658 84044 -1594
rect 69804 -4036 69860 -3972
rect 70081 -4036 70102 -3972
rect 83551 -4036 84044 -3972
rect 58988 -4160 58989 -4096
rect 59053 -4160 59054 -4096
rect 83379 -6516 83380 -6452
rect 83444 -6516 83445 -6452
rect 58306 -6640 58866 -6576
rect 58930 -6640 58989 -6576
rect 83454 -8996 83503 -8932
rect 83567 -8996 84023 -8932
rect 58988 -9120 58989 -9056
rect 59053 -9120 59054 -9056
rect 83379 -11476 83380 -11412
rect 83444 -11476 83445 -11412
rect 83551 -11600 83626 -11536
rect 83690 -11600 83700 -11536
rect 58383 -13956 58879 -13892
rect 83502 -14080 83503 -14016
rect 83567 -14080 83568 -14016
rect 58346 -16436 58879 -16372
rect 60425 -16416 60485 -16155
rect 83551 -16436 83626 -16372
rect 83690 -16436 84056 -16372
rect 83379 -16560 83380 -16496
rect 83444 -16560 83445 -16496
rect 58988 -18916 58989 -18852
rect 59053 -18916 59054 -18852
rect 58865 -21396 58866 -21332
rect 58930 -21396 58931 -21332
rect 83379 -21520 83380 -21456
rect 83444 -21520 83445 -21456
rect 83514 -21520 84033 -21456
rect 58243 -23876 58911 -23812
rect 83610 -24000 84044 -23936
<< via3 >>
rect 83379 18182 83445 18246
rect 58988 15826 59052 15890
rect 83504 15702 83568 15766
rect 58866 13346 58930 13410
rect 83379 13222 83445 13286
rect 58989 10866 59053 10930
rect 58743 10742 58807 10806
rect 72347 10742 72565 10806
rect 58866 8386 58930 8450
rect 58743 5906 58807 5970
rect 58989 5782 59053 5846
rect 83379 3426 83445 3490
rect 58866 3302 58930 3366
rect 83504 946 83568 1010
rect 58989 822 59053 886
rect 83379 -1534 83445 -1470
rect 69860 -1658 70081 -1594
rect 69860 -4036 70081 -3972
rect 58989 -4160 59053 -4096
rect 83380 -6516 83444 -6452
rect 58866 -6640 58930 -6576
rect 83503 -8996 83567 -8932
rect 58989 -9120 59053 -9056
rect 83380 -11476 83444 -11412
rect 83626 -11600 83690 -11536
rect 83503 -14080 83567 -14016
rect 83626 -16436 83690 -16372
rect 83380 -16560 83444 -16496
rect 58989 -18916 59053 -18852
rect 83503 -19040 83567 -18976
rect 58866 -21396 58930 -21332
rect 83380 -21520 83444 -21456
rect 58989 -23876 59053 -23812
<< metal4 >>
rect 83382 18247 83442 18387
rect 83378 18246 83446 18247
rect 83378 18182 83379 18246
rect 83445 18182 83446 18246
rect 83378 18181 83446 18182
rect 58991 15891 59051 15924
rect 58987 15890 59053 15891
rect 58987 15826 58988 15890
rect 59052 15826 59053 15890
rect 58987 15825 59053 15826
rect 58868 13411 58928 13458
rect 58865 13410 58931 13411
rect 58865 13346 58866 13410
rect 58930 13346 58931 13410
rect 58865 13345 58931 13346
rect 58745 10807 58805 10818
rect 58742 10806 58808 10807
rect 58742 10742 58743 10806
rect 58807 10742 58808 10806
rect 58742 10741 58808 10742
rect 58745 5971 58805 10741
rect 58868 8451 58928 13345
rect 58991 10931 59051 15825
rect 83382 13287 83442 18181
rect 83506 15767 83566 15787
rect 83503 15766 83569 15767
rect 83503 15702 83504 15766
rect 83568 15702 83569 15766
rect 83503 15701 83569 15702
rect 83378 13286 83446 13287
rect 83378 13222 83379 13286
rect 83445 13222 83446 13286
rect 83378 13221 83446 13222
rect 58988 10930 59054 10931
rect 58988 10866 58989 10930
rect 59053 10866 59054 10930
rect 58988 10865 59054 10866
rect 58865 8450 58931 8451
rect 58865 8386 58866 8450
rect 58930 8386 58931 8450
rect 58865 8385 58931 8386
rect 58742 5970 58808 5971
rect 58742 5906 58743 5970
rect 58807 5906 58808 5970
rect 58742 5905 58808 5906
rect 58745 5873 58805 5905
rect 58868 3367 58928 8385
rect 58991 5847 59051 10865
rect 72346 10806 72566 10807
rect 72346 10742 72347 10806
rect 72565 10742 72566 10806
rect 72346 10741 72566 10742
rect 72425 10476 72485 10741
rect 58988 5846 59054 5847
rect 58988 5782 58989 5846
rect 59053 5782 59054 5846
rect 58988 5781 59054 5782
rect 58865 3366 58931 3367
rect 58865 3302 58866 3366
rect 58930 3302 58931 3366
rect 58865 3301 58931 3302
rect 58868 3274 58928 3301
rect 58991 887 59051 5781
rect 83382 3491 83442 13221
rect 83378 3490 83446 3491
rect 83378 3426 83379 3490
rect 83445 3426 83446 3490
rect 83378 3425 83446 3426
rect 58988 886 59054 887
rect 58988 822 58989 886
rect 59053 822 59054 886
rect 58988 821 59054 822
rect 58991 792 59051 821
rect 60025 -1924 60085 -1204
rect 69945 -1593 70005 -1144
rect 69859 -1594 70082 -1593
rect 69859 -1658 69860 -1594
rect 70081 -1658 70082 -1594
rect 69859 -1659 70082 -1658
rect 82345 -1924 82405 -1204
rect 83382 -1469 83442 3425
rect 83506 1011 83566 15701
rect 83503 1010 83569 1011
rect 83503 946 83504 1010
rect 83568 946 83569 1010
rect 83503 945 83569 946
rect 83506 935 83566 945
rect 83378 -1470 83446 -1469
rect 83378 -1534 83379 -1470
rect 83445 -1534 83446 -1470
rect 83378 -1535 83446 -1534
rect 83382 -1558 83442 -1535
rect 60935 -2845 61655 -2785
rect 63415 -2845 64135 -2785
rect 65895 -2845 66615 -2785
rect 73335 -2845 74055 -2785
rect 75815 -2845 76535 -2785
rect 78295 -2845 79015 -2785
rect 80775 -2845 81495 -2785
rect 58991 -4095 59051 -4071
rect 58988 -4096 59054 -4095
rect 58988 -4160 58989 -4096
rect 59053 -4160 59054 -4096
rect 58988 -4161 59054 -4160
rect 58868 -6575 58928 -6540
rect 58865 -6576 58931 -6575
rect 58865 -6640 58866 -6576
rect 58930 -6640 58931 -6576
rect 58865 -6641 58931 -6640
rect 58868 -21331 58928 -6641
rect 58991 -9055 59051 -4161
rect 60025 -4426 60085 -3706
rect 69945 -3971 70005 -3705
rect 69859 -3972 70082 -3971
rect 69859 -4036 69860 -3972
rect 70081 -4036 70082 -3972
rect 69859 -4037 70082 -4036
rect 69945 -4426 70005 -4037
rect 82345 -4426 82405 -3706
rect 83382 -6451 83442 -6402
rect 83379 -6452 83445 -6451
rect 83379 -6516 83380 -6452
rect 83444 -6516 83445 -6452
rect 83379 -6517 83445 -6516
rect 58988 -9056 59054 -9055
rect 58988 -9120 58989 -9056
rect 59053 -9120 59054 -9056
rect 58988 -9121 59054 -9120
rect 58991 -18851 59051 -9121
rect 83382 -11411 83442 -6517
rect 83505 -8931 83565 -8920
rect 83502 -8932 83568 -8931
rect 83502 -8996 83503 -8932
rect 83567 -8996 83568 -8932
rect 83502 -8997 83568 -8996
rect 83379 -11412 83445 -11411
rect 83379 -11476 83380 -11412
rect 83444 -11476 83445 -11412
rect 83379 -11477 83445 -11476
rect 69945 -14346 70005 -13626
rect 68375 -15256 69095 -15196
rect 70855 -15256 71575 -15196
rect 69945 -16826 70005 -16106
rect 83382 -16495 83442 -11477
rect 83505 -14015 83565 -8997
rect 83628 -11535 83688 -11501
rect 83625 -11536 83691 -11535
rect 83625 -11600 83626 -11536
rect 83690 -11600 83691 -11536
rect 83625 -11601 83691 -11600
rect 83502 -14016 83568 -14015
rect 83502 -14080 83503 -14016
rect 83567 -14080 83568 -14016
rect 83502 -14081 83568 -14080
rect 83379 -16496 83445 -16495
rect 83379 -16560 83380 -16496
rect 83444 -16560 83445 -16496
rect 83379 -16561 83445 -16560
rect 58988 -18852 59054 -18851
rect 58988 -18916 58989 -18852
rect 59053 -18916 59054 -18852
rect 58988 -18917 59054 -18916
rect 58865 -21332 58931 -21331
rect 58865 -21396 58866 -21332
rect 58930 -21396 58931 -21332
rect 58865 -21397 58931 -21396
rect 58868 -21567 58928 -21397
rect 58991 -23811 59051 -18917
rect 83382 -21455 83442 -16561
rect 83505 -18975 83565 -14081
rect 83628 -16371 83688 -11601
rect 83625 -16372 83691 -16371
rect 83625 -16436 83626 -16372
rect 83690 -16436 83691 -16372
rect 83625 -16437 83691 -16436
rect 83628 -16455 83688 -16437
rect 83502 -18976 83568 -18975
rect 83502 -19040 83503 -18976
rect 83567 -19040 83568 -18976
rect 83502 -19041 83568 -19040
rect 83505 -19066 83565 -19041
rect 83379 -21456 83445 -21455
rect 83379 -21520 83380 -21456
rect 83444 -21520 83445 -21456
rect 83379 -21521 83445 -21520
rect 83382 -21539 83442 -21521
rect 58988 -23812 59054 -23811
rect 58988 -23876 58989 -23812
rect 59053 -23876 59054 -23812
rect 58988 -23877 59054 -23876
rect 58991 -24043 59051 -23877
use cap_array_half  cap_array_half_0
timestamp 1718210529
transform -1 0 164043 0 -1 -5781
box 80293 -26673 105363 -4081
use cap_array_half  cap_array_half_1
timestamp 1718210529
transform 1 0 -21613 0 1 151
box 80293 -26673 105363 -4081
use caparray_connect_near  caparray_connect_near_0
timestamp 1717937330
transform -1 0 151643 0 -1 -28101
box 80427 -26673 82908 -26177
use cdac_cross2_short  cdac_cross2_short_0
timestamp 1718207857
transform 1 0 14880 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_1
timestamp 1718207857
transform 1 0 -4960 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_2
timestamp 1718207857
transform 1 0 -2480 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_3
timestamp 1718207857
transform 1 0 0 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_6
timestamp 1718207857
transform 1 0 7440 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_7
timestamp 1718207857
transform 1 0 9920 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_8
timestamp 1718207857
transform 1 0 12400 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross_short  cdac_cross_short_0
timestamp 1718207857
transform 0 1 62881 -1 0 64691
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_1
timestamp 1718207857
transform 1 0 14880 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_2
timestamp 1718207857
transform 1 0 -4960 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_3
timestamp 1718207857
transform 1 0 -2480 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_4
timestamp 1718207857
transform 1 0 0 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_5
timestamp 1718207857
transform 1 0 2480 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_6
timestamp 1718207857
transform 1 0 4960 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_7
timestamp 1718207857
transform 1 0 7440 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_8
timestamp 1718207857
transform 1 0 9920 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_9
timestamp 1718207857
transform 1 0 12400 0 1 -22320
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_10
timestamp 1718207857
transform 0 -1 57229 1 0 -75281
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_11
timestamp 1718207857
transform 0 -1 57229 1 0 -77761
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_12
timestamp 1718207857
transform 0 -1 57229 1 0 -87681
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_13
timestamp 1718207857
transform 0 -1 57229 1 0 -82721
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_14
timestamp 1718207857
transform 0 -1 57229 1 0 -85201
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_15
timestamp 1718207857
transform 0 1 62881 -1 0 82051
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_16
timestamp 1718207857
transform 0 1 85201 -1 0 82051
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_17
timestamp 1718207857
transform 0 1 85201 -1 0 47309
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_18
timestamp 1718207857
transform 0 1 85201 -1 0 49789
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_19
timestamp 1718207857
transform 0 1 85201 -1 0 52269
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_20
timestamp 1718207857
transform 0 1 85201 -1 0 54749
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_21
timestamp 1718207857
transform 0 1 85201 -1 0 57229
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_22
timestamp 1718207857
transform 0 1 85201 -1 0 59709
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_23
timestamp 1718207857
transform 0 1 85201 -1 0 62189
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_24
timestamp 1718207857
transform 0 1 85201 -1 0 64691
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_25
timestamp 1718207857
transform 0 1 85201 -1 0 67171
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_26
timestamp 1718207857
transform 0 1 85201 -1 0 69651
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_27
timestamp 1718207857
transform 0 1 85201 -1 0 72131
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_28
timestamp 1718207857
transform 0 1 85201 -1 0 74611
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_29
timestamp 1718207857
transform 0 1 85201 -1 0 77091
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_30
timestamp 1718207857
transform 0 1 85201 -1 0 79571
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_31
timestamp 1718207857
transform 0 1 85201 -1 0 44829
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_32
timestamp 1718207857
transform 0 -1 57229 1 0 -80241
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_33
timestamp 1718207857
transform 0 -1 57229 1 0 -72801
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_34
timestamp 1718207857
transform 0 -1 57229 1 0 -70321
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_35
timestamp 1718207857
transform 0 1 62881 -1 0 72131
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_36
timestamp 1718207857
transform 0 1 62881 -1 0 69651
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_37
timestamp 1718207857
transform 0 1 62881 -1 0 67171
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_38
timestamp 1718207857
transform 0 1 62881 -1 0 79571
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_39
timestamp 1718207857
transform 0 1 62881 -1 0 77091
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_40
timestamp 1718207857
transform 0 1 62881 -1 0 74611
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_41
timestamp 1718207857
transform 1 0 14880 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_42
timestamp 1718207857
transform 1 0 12400 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_43
timestamp 1718207857
transform 1 0 9920 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_44
timestamp 1718207857
transform 1 0 7440 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_45
timestamp 1718207857
transform 1 0 4960 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_46
timestamp 1718207857
transform 1 0 2480 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_47
timestamp 1718207857
transform 1 0 0 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_48
timestamp 1718207857
transform 1 0 -2480 0 1 22342
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_49
timestamp 1718207857
transform 1 0 -4960 0 1 22342
box 65895 -3386 66615 -2266
use cdac_ratioed_cap  cdac_ratioed_cap_0
array 0 9 2480 0 0 2797
timestamp 1717944067
transform 1 0 -21716 0 1 29649
box 80396 -33851 83146 -31078
<< labels >>
flabel comment 83579 -11569 83579 -11569 0 FreeSans 800 0 0 0 D1
flabel comment 58853 -21366 58853 -21366 0 FreeSans 800 0 0 0 D2
flabel comment 58858 -6610 58858 -6610 0 FreeSans 800 0 0 0 D2
flabel comment 83585 -19010 83585 -19010 0 FreeSans 800 0 0 0 D3
flabel comment 83587 -14052 83587 -14052 0 FreeSans 800 0 0 0 D3
flabel comment 83582 -8968 83582 -8968 0 FreeSans 800 0 0 0 D3
flabel comment 58850 -23849 58850 -23849 0 FreeSans 800 0 0 0 D4
flabel comment 58864 -18883 58864 -18883 0 FreeSans 800 0 0 0 D4
flabel comment 58859 -9083 58859 -9083 0 FreeSans 800 0 0 0 D4
flabel comment 58859 -4132 58859 -4132 0 FreeSans 800 0 0 0 D4
flabel comment 83577 -21482 83577 -21482 0 FreeSans 800 0 0 0 D5
flabel comment 83566 -16524 83566 -16524 0 FreeSans 800 0 0 0 D5
flabel comment 83566 -11441 83566 -11441 0 FreeSans 800 0 0 0 D5
flabel comment 83566 -6489 83566 -6489 0 FreeSans 800 0 0 0 D5
flabel comment 83583 10775 83583 10775 0 FreeSans 800 0 0 0 VSS
flabel comment 58847 5934 58847 5934 0 FreeSans 800 0 0 0 D7
flabel comment 58847 10766 58847 10766 0 FreeSans 800 0 0 0 D7
flabel comment 83575 8295 83575 8295 0 FreeSans 800 0 0 0 D6
flabel comment 83587 977 83587 977 0 FreeSans 800 0 0 0 D8
flabel comment 83576 15736 83576 15736 0 FreeSans 800 0 0 0 D8
flabel comment 58837 3322 58837 3322 0 FreeSans 800 0 0 0 D9
flabel comment 58843 8414 58843 8414 0 FreeSans 800 0 0 0 D9
flabel comment 58859 13375 58859 13375 0 FreeSans 800 0 0 0 D9
flabel comment 83588 -1497 83588 -1497 0 FreeSans 800 0 0 0 D10
flabel comment 83571 13253 83571 13253 0 FreeSans 800 0 0 0 D10
flabel comment 83575 18212 83575 18212 0 FreeSans 800 0 0 0 D10
flabel comment 58855 851 58855 851 0 FreeSans 800 0 0 0 D11
flabel comment 58855 5813 58855 5813 0 FreeSans 800 0 0 0 D11
flabel comment 58855 10892 58855 10892 0 FreeSans 800 0 0 0 D11
flabel comment 58859 15862 58859 15862 0 FreeSans 800 0 0 0 D11
flabel comment 58877 -13922 58877 -13922 0 FreeSans 800 0 0 0 D0
flabel comment 58889 -16402 58889 -16402 0 FreeSans 800 0 0 0 VSS
flabel comment 58868 -11570 58868 -11570 0 FreeSans 800 0 0 0 D1
flabel comment 83547 -16401 83547 -16401 0 FreeSans 800 0 0 0 D1
flabel comment 83564 3460 83564 3460 0 FreeSans 800 0 0 0 D10
flabel metal3 58344 10742 58544 10806 0 FreeSans 480 0 0 0 D7
port 11 nsew
flabel metal3 58258 3302 58458 3366 0 FreeSans 480 0 0 0 D9
port 4 nsew
flabel metal3 58324 15826 58516 15890 0 FreeSans 480 0 0 0 D11
port 14 nsew
flabel metal3 58308 -6640 58508 -6576 0 FreeSans 480 0 0 0 D2
port 8 nsew
flabel metal3 58386 -13956 58545 -13892 0 FreeSans 480 0 0 0 D0
port 1 nsew
flabel metal3 58244 -23876 58444 -23812 0 FreeSans 480 0 0 0 D4
port 2 nsew
flabel metal3 83830 -21520 84030 -21456 0 FreeSans 480 0 0 0 D5
port 5 nsew
flabel metal3 83854 -16436 84054 -16372 0 FreeSans 480 0 0 0 D1
port 6 nsew
flabel metal3 83822 -8996 84022 -8932 0 FreeSans 480 0 0 0 D3
port 12 nsew
flabel metal3 83840 -4036 84040 -3972 0 FreeSans 480 0 0 0 VP1
port 3 nsew
flabel metal3 83848 -1658 84044 -1594 0 FreeSans 480 0 0 0 VP2
port 7 nsew
flabel metal3 83780 946 83980 1010 0 FreeSans 480 0 0 0 D8
port 0 nsew
flabel metal3 83798 8262 83997 8326 0 FreeSans 480 0 0 0 D6
port 9 nsew
flabel metal3 58348 -16436 58545 -16372 0 FreeSans 480 0 0 0 VSS
port 10 nsew
flabel metal3 83928 18182 84120 18246 0 FreeSans 480 0 0 0 D10
port 13 nsew
<< end >>
