** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/sky130_ef_ip__cdac10bit.sch
.subckt sky130_ef_ip__cdac10bit SELD0 SELD1 SELD2 SELD3 SELD4 SELD5 SELD6 SELD7 SELD8 SELD9 VDD DVDD DVSS VSS VH VL OUT RST EN
*.PININFO SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VDD:B DVDD:B DVSS:B VH:B VL:B VSS:B
*+ RST:I EN:I OUT:O
x4 D8 D0 D4 VP1 D9 D5 D1 VP2 D2 D6 VSS D7 D3 EF_BANK_CAP_10
x3 D0 SELD0 D1 SELD1 SELD2 D2 SELD3 SELD4 D3 SELD5 D4 SELD6 SELD7 D5 SELD8 D6 SELD9 D7 D8 D9 VDD DVDD DVSS VH VL VSS
+ EF_AMUX0201_ARRAY1
x1 VP1 VP2 VDD DVDD VSS RST DVSS EF_SW_RST
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=24
x5 VDD OUT EN3V VSS VP2 DVSS follower_amp
XC1 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=24
x2 EN DVDD DVSS DVSS VDD VDD EN3V sky130_fd_sc_hvl__lsbuflv2hv_1
.ends

* expanding   symbol:  EF_BANK_CAP_10.sym # of pins=13
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_BANK_CAP_10.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_BANK_CAP_10.sch
.subckt EF_BANK_CAP_10 D8 D0 D4 VP1 D9 D5 D1 VP2 D2 D6 VSS D7 D3
*.PININFO D0:B D1:B D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B VSS:B VP1:B VP2:B
x4 VP1 VSS D0 D1 D2 D3 D4 EF_LSB_CAP
x1 D8 D5 D9 VP2 D6 VSS D7 EF_MSB_CAP
x2 VP1 VP2 VSS EF_SC_CAP
.ends


* expanding   symbol:  EF_AMUX0201_ARRAY1.sym # of pins=26
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_AMUX0201_ARRAY1.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_AMUX0201_ARRAY1.sch
.subckt EF_AMUX0201_ARRAY1 D0 SELD0 D1 SELD1 SELD2 D2 SELD3 SELD4 D3 SELD5 D4 SELD6 SELD7 D5 SELD8 D6 SELD9 D7 D8 D9 VDD DVDD DVSS
+ VH VL VSS
*.PININFO VDD:B DVDD:B DVSS:B VH:B VL:B SELD0:I SELD1:I SELD2:I SELD3:I SELD4:I SELD5:I SELD6:I SELD7:I SELD8:I SELD9:I VSS:B D0:B
*+ D1:B D2:B D3:B D4:B D5:B D6:B D7:B D8:B D9:B
x2 VDD DVDD D0 VSS VH VL SELD0 DVSS EF_AMUX21x
x1 VDD DVDD D1 VSS VH VL SELD1 DVSS EF_AMUX21x
x3 VDD DVDD D2 VSS VH VL SELD2 DVSS EF_AMUX21x
x4 VDD DVDD D3 VSS VH VL SELD3 DVSS EF_AMUX21x
x5 VDD DVDD D4 VSS VH VL SELD4 DVSS EF_AMUX21x
x8 VDD DVDD D5 VSS VH VL SELD5 DVSS EF_AMUX21x
x9 VDD DVDD D6 VSS VH VL SELD6 DVSS EF_AMUX21x
x10 VDD DVDD D7 VSS VH VL SELD7 DVSS EF_AMUX21x
x11 VDD DVDD D8 VSS VH VL SELD8 DVSS EF_AMUX21x
x12 VDD DVDD D9 VSS VH VL SELD9 DVSS EF_AMUX21x
.ends


* expanding   symbol:  EF_SW_RST.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_SW_RST.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_SW_RST.sch
.subckt EF_SW_RST VP1 VP2 AVDD DVDD AVSS RST DVSS
*.PININFO AVSS:B DVDD:B AVDD:B VP1:B VP2:B RST:I DVSS:B
x1 AVSS RST VP2 AVSS AVDD DVDD DVSS simple_analog_switch_ena1v8
x2 AVSS RST VP1 AVSS AVDD DVDD DVSS simple_analog_switch_ena1v8
.ends


* expanding   symbol:  ../dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sym # of pins=6
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sch
.subckt follower_amp vdd out ena vss in vsub
*.PININFO in:I vdd:I vss:I out:O ena:I vsub:I
XM4 pdrv1 net1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM5 vdd net1 net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM10 vss nbias nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=4 m=1
XM20 out pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=280 nf=280 m=1
XM22 out ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=4 m=1
XM24 pbias nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM25 vdd pbias pbias vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM26 vcomp pbias vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM27 net2 out vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM28 vcomp in ndrv vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM29 ndrv net2 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM30 vss net2 net2 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM1 net1 out vcomn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 vcomn1 in pdrv1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 pdrv2 net3 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM6 vdd net3 net3 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM7 vcomn2 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM12 vdd pdrv2 out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=20 m=1
XXD1 vss in sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=4e6
XM13 net4 ena nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XXD2 vss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=4e6
XM11 pdrv2 in vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM9 net3 out vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM8 vcomn1 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR2 net4 vdd vss sky130_fd_pr__res_xhigh_po_0p35 L=35 mult=1 m=1
.ends


* expanding   symbol:  EF_LSB_CAP.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_LSB_CAP.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_LSB_CAP.sch
.subckt EF_LSB_CAP VP1 VSS D0 D1 D2 D3 D4
*.PININFO VP1:B D0:B D1:B D2:B D3:B D4:B VSS:B
XC1 VP1 VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC2 VP1 D0 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC8 VSS VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VP1 D1 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC4 VP1 D2 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC5 VP1 D3 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC7 VP1 D4 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC9 D0 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC10 D1 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC11 D2 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC12 D3 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC13 D4 VP1 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC14 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
.ends


* expanding   symbol:  EF_MSB_CAP.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_MSB_CAP.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_MSB_CAP.sch
.subckt EF_MSB_CAP D8 D5 D9 VP2 D6 VSS D7
*.PININFO D5:B D6:B D7:B D8:B D9:B VP2:B VSS:B
XC1 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC2 D5 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC3 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=32
XC4 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=32
XC5 VSS VSS sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=1
XC6 VP2 D5 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=1
XC7 VP2 D6 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=2
XC8 VP2 D7 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=4
XC9 VP2 D8 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=8
XC10 VP2 D9 sky130_fd_pr__cap_mim_m3_1 W=7 L=7 m=16
XC11 D6 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=2
XC12 D7 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=4
XC13 D8 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=8
XC14 D9 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7 m=16
.ends


* expanding   symbol:  EF_SC_CAP.sym # of pins=3
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_SC_CAP.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_SC_CAP.sch
.subckt EF_SC_CAP VP1 VP2 VSS
*.PININFO VP1:B VP2:B VSS:B
XC13 VP2 VP1 sky130_fd_pr__cap_mim_m3_1 W=7 L=7.225 m=1
XC6 VSS VSS sky130_fd_pr__cap_mim_m3_1 W=7 L=7.225 m=7
XC1 net1 net2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7.225 m=1
XC2 VP1 VP2 sky130_fd_pr__cap_mim_m3_2 W=7 L=7.225 m=1
.ends


* expanding   symbol:  EF_AMUX21x.sym # of pins=8
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_AMUX21x.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/xschem/EF_AMUX21x.sch
.subckt EF_AMUX21x vdd3p3 vdd1p8 vo vss a b sel dvss
*.PININFO sel:I vo:B vdd3p3:B vss:B vdd1p8:B dvss:B a:B b:B
x1 vss sel vo a vdd3p3 vdd1p8 dvss simple_analog_switch_ena1v8
x4 vss selp vo b vdd3p3 vdd1p8 dvss simple_analog_switch_ena1v8
x5 sel vss vss vdd1p8 vdd1p8 selp sky130_fd_sc_hvl__inv_2
.ends


* expanding   symbol:  ../dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sym
** sch_path: /home/tim/gits/sky130_ef_ip__cdac3v_10bit/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sch
.subckt simple_analog_switch_ena1v8 avss on out in avdd dvdd dvss
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B
x2 on dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
XD1 dvss on sky130_fd_pr__diode_pw2nd_05v5 area=2.304e11 perim=1.92e6
x3 net1 net2 avss out in avdd simple_analog_switch
x1 net3 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x4 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
.ends


* expanding   symbol:  simple_analog_switch.sym # of pins=6
** sym_path: /home/tim/gits/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sym
** sch_path: /home/tim/gits/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sch
.subckt simple_analog_switch on off vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B off:I
XM1 in on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 in off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=4 m=1
XM3 out off out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 out on out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM5 in off in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 in on in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
.ends

.end
