magic
tech sky130A
magscale 1 2
timestamp 1718225130
<< error_p >>
rect 81108 -26399 81428 -26353
rect 81108 -26635 81150 -26399
rect 81108 -26673 81428 -26635
<< metal3 >>
rect 82038 -26443 82098 -26177
rect 80427 -26507 81151 -26443
rect 81385 -26507 82908 -26443
rect 80427 -26631 82908 -26567
<< via3 >>
rect 81151 -26507 81385 -26443
<< via4 >>
rect 81150 -26443 81386 -26399
rect 81150 -26507 81151 -26443
rect 81151 -26507 81385 -26443
rect 81385 -26507 81386 -26443
rect 81150 -26635 81386 -26507
<< metal5 >>
rect 81108 -26399 81428 -26354
rect 81108 -26635 81150 -26399
rect 81386 -26635 81428 -26399
rect 81108 -26673 81428 -26635
<< end >>
